// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:35 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
T8vGdZUSUQZDWoFL7Jrs7qJpDxMlLMtVSX3QxgKap1kudbeB+hz2SzrxuykvHxaN
NruBFUrlcgox0nBfPMh03bAILgo/mPBtofzEMNatKvcru0FUF6dFD7DfLdolDb4d
xTyLug63qVFWzLFNUL9NnglCmuMXtslks+53C07FTrk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35392)
RseSsVzThaXC9acVswduNBgOfqcZoynGbsjDz4SYy9XMEkJL1GfCCaYGnVOWvBR7
0cIs16WFhNOis0KCfQfGw6SZPVrUsFIhz6Z0L+wrw6xYg05NciHWAXuvEBHyb2N+
pRIEUd6oul6lUccjnlSYU3231CI/xMf4IFLD1Wq8bNXJwCVbaaZ+20T3EKmHb9tu
jPq+QfZzPvxx8joRtWVibCfx2uSVej9IincDFTEdaAREuI3S3//IYCV68lXM0o9u
dtucm5nfXaZyF9vkYvFeW/l/2Ij4CmGQ7uu3uYGdJ5fnhntQqpxi/vpLhvpn2XdC
vwnhewNkYLb3nHcFiWlICSaNEDzdH7sl/uFIbn0kPdUi9pXTDgSeVttov8VfVlj6
UualfTkrXVHwwn2s89VtxucOVGCcwiB2qLecHqQD5Ae1IJKMA/luqGIAE12nJk+s
lnJWLJ3J0UMpSi5SwsYVGC5M0Ds2nUVhPt8E6VvlCse2Gpyu4g4ySd0hmxZ/pUKw
9MQfx94393XrADrYSavMxYKEMFqUHNEaaRGR4AUFKCi8tlSxKuarObu6a9zOwOaE
OpV8GBAwguTEl3vYboZdrnhY2SNqja+V7cncJhfsPscT12IPfXvXuBkGEtshQZ07
+kilURv6gx4JADyTsjQPRyW9N/oOIBF88H1oj8ZogmA2GeXjBAVA2zJKWXe3Gi0c
mL8+dvb9lv5T4RUvPi1F6R/VdGAp8Mqq8fueDM/INNPgMGQbiXoQmviALgVxm9js
29QrspeLzlKw6o11QiSUVf2Zaz7VNzij5cV7nbnZS78B3RpzNWC3cJrIL6+nPoDt
2Nlz+8kFslYL+M9K7izTz2VrpCU30A/7ozvWNsIQzSONGlY+5V1qsu1/ntpnChiG
hs5/Du5XErlgSVgosQL7X/GqCohDOonyoRy9NwKKlvwjYBxKK1rm8bZwyCPLnQnd
STBC5Z6Q953xMq8LL+L+XFJJifxRis1J693tSyiFPraOSHcvOdQZzkfWgrY/GoYf
rl4q65MX+uOlzyuqmuOcAcSU2dP2fmSbY0C2aewlD5M/frLDFcJuzfGI+4ZqD9RF
ShIgAn1goOAQOHfTyLFioYXs3s6YsRIiAHDtH7pjCpHczjvaXtjy+iXSgofhfO+g
KPvPyStZdYJM1rhnlLcj2r0BZ3s6haGmU34GC9YyesjuHBNbHnBcAy94Nb2y6u7J
AH+HBAHyNR9vj7WOjdfOUOPdh4I+y6VacNpElvkAMWjKjNUGO9QLshU7Px7aSPB2
DnhmLLK1Q0GqzvylE+A7jgAGsbjomdP4YmYcAwhZYAN9f3F8TDC0M5/QkeC8pASv
06CjnunbG8VjdXf+IocItLpaJOILWQwS4dv08LDFItJ9ps9bHnZRKKnrv84rA+nu
qBSkwdCKPWmgFE9RBnb4puV9/lp2O/VFJY4yo+Tz65E36zjIPDiMAYwCfS737FJr
K1TJrahPfnwhFQlWje6LXRoE39dPOhPCbPAfFgj6lCbSzWOnnz7j9PvcxL6fy48P
JmJFYJbi4SI2YeKaQws5TguEZEU0ncTP1M4aoBJ1jkD4oYywooowpHWa0N5wcNWo
LIzVE1G0aipfRSON1m+tA3r40Ul9mzHxuY6069tg70CV3FA+2iDpaUKFBt5EMige
2Wt6zDTxRXFe2aGp+Ydvg0gS513pPl8psyAOL2nulQNR+0CB9rmLgsY9zoVkmI36
WiLSbYBcceVN7tw7BlT/NgckGdo9OqyaSFLD9NS2epVytxQxAHRoACkNnESllJty
r2PFx3zsWNokoaH+66nZlt4RwDW+vZLeAbkyVy3Cja1LpJwvxBfR6eFLXE1Txfvr
2jjE8cZzqdukTo4K46e4ZN4dRa8H0TtGjfh6Q5EKXaqQGRywj+PcTmUyB5dDXmWo
SXZWkPLIb5jD20E9f41hLOmut68P78xLRQDRYCmitkaae7oLOA60rKDdMwYntEaD
Xwd1Jomq1hhOFoiDKnfSYDcM5KBfj7e310Q2zU3f7RDI4e9bVXAMISABVdcdK5As
qB4+RQw4kLLONVyg9fOfftgJa/wUKQ3ucfvK5gZfIH6acv9bYRDfykivH4duxu+B
tKTNFelJbw7GfOb3YGLioJ6TunsmKl8FJvm1NZWTG+heN/vpsquhIu59M4aSNDm1
ni8NSGVS6bIq4POYC6FUMFkjWi5nR7Q8y0nA5a4gBrh2Ws3UK60Ue6k9V9QEzQSR
14BrYV6ySkrBf6MeYzxZ8/iUzSN5g33sBtZJUurl8a8ns7PpewLwpRt+indhdx/4
Wz+Lb5xU5VfItDwkVtZ770Acn4y3O4kylRNIhzFIi9184AWPIqpXTviKQ18kohAd
B5hcy5h4yZrL2SWwkxS3sJX368LK57FQ91NEi/PTXLB5aQ17BNaS+gF0Wn3RxKS+
HJvBUi1puBbLU5ldKicsCd/iN6WLGQE5f6+8VlixAah6OjfOAVHVuXZEQiLArVIE
WB+9CaUuwN7bcCED/C8FlFy/Z/K+541Ahnp/oNMjiwwogz6zvlITeiSqG7wGbjPK
sNSolYyGhVniRZDlAeioBjdjGrYnUt70416jq5Tf2beyN5NQnawkq3Ivw47nihFB
T//qa7Oh4SkLr0HWxpg7ouoH4gwhOQwG3ePbYGdO+yGssFzh7MVqG7RzHL2YS5mM
J5+CAQ9ktShPW6/akjwhzpIIVrGkjEwK4qgzUBLjoYMVuqeTQXr1+uwGZQkB5mug
TzJR0rlanxvHzs/T8EDF14Fc0DuF1wC4tUcENIqWREJCOrEsapWxhGkNgd+C1beW
Yw7z7zBW93huBH51a1wckp6ShI1r4YEVQEjY6Dmjt5VWOKd0baDSB0TgvdpYxzgw
D46+H7LAIamtotXR9hwhL9l3rc1yjIQXVfWc8kMAK/R8ywSsVPXoBt4j6vKQstlf
PKr87iJTw6X9pWrdd2sJobFketSehHFaEx6wl7lkMuADpCrU6K+F7dIZHoQdSdFX
+UkvUQEUvPBI9PWoDP69PsaLmd9mGJ9caT3w3AjqTYShqHEEnXEnJvSc7UbCzajz
9JITGWk1aNpCsK0sJdQHbEX/V1STuL+Fy4gL7tGBKE8UYVhJnaf4gQKvSvOuvUh8
nEbd3NrDuGn0LIPA4DrSpYe5YeVAf0mhidswkNhjaIYItM4kxiIl3r9bGRMQ6QMg
2lIIdZVRNpemT6Uo7ZWRg1u7nkaXv3IbQSk89oSa15cUl6JSiHKw6xsFR1kNww5s
2U/C61R7hk4A6kHVrPntUNwQwRRma4/fxt0TK0v3+VJqmeMtD7GWHktyl3mnFxr4
okQGTMuMc6HnxxF9eVQGa99TpqyvTU3venwo2+D4YN/UwfH4o3lG7ZH8UC+GXS36
D8hQ6M+2koDaHs+bdndvXbVG3hLw76GYQoEuYEJYxHI0ihV2mrbWj44otx9h6U57
a7eBgtsrux0soefR40kYaHHM8zTr/GYuy6EYo5zlJfgEQUOz6W7/H3BZE87mPGiR
yp5eKoHfLs/sH0wv3DY55viNF8u3Ur6QhpyGZGk9dGjtqqDC6oSRX9YEYHI94rYT
1QkFKcksQqd8YIsIWLh0XWoZVlCni/ftqv1CiiZnLvoARGkyk60LfmT+fqg0iIeP
9dLuvExd+FKOOzyH6/+/90NPdP4WYsQUxj0/IguUq8TspMkKK/91e8xFgNlYzFjY
vzYpaIbGmfj4y/Wg99J1c5qKpWca3QpOhDXdt4Gswlf7bD7GMa20kkEABYpt0j7y
sSK9sO24bnZJ3ym+gwE+WLqO5UXgVzdkqE071CLp9wdlPxh21IxpGyDjWqsL2K04
AkYL5Cpd1dT/IS0P+PmcjmlNXpmyz5hJrkeiar7ozyYpLto2pkMAkGJodJNFOOfa
8nB77nG/eKVqbYot3ecRPJ4Q2H+UKWipcAJjCVYgkVA1jCaAeLddrL3BhmOR4v9F
54Ps2ocUGh+SPHWepKT3F/wG96d8ddzPL5jo1n44AiYSmU8TEJMfQV4T/n2QMZfy
zyZx06WWYBD6/b7QjLhqWJqEOmuk+Vm0V/Mhk/kwJ767Inm8tP+tY3jE8PFPq2qE
Yt08/XanuAHFo54jrWzMBpyB0o+99S8JS0mhhuuv6815tltO935c3DFvUsB7ONr4
IyRs08j1BbIHSsQ6lFaNCm/c2WYbGQE6mcmwtRGCs72vOnVnJPNaRXNNTH9hXn7O
r5klaujeG/bb0TgElH2uLIyqL4GTp37iSvbWAR99nFi1N4TLziaZd7SW2RvGQfux
HZ7FrKlWDSjFWAbd0Rvzu9nyzuU0p4SbDLs+tWF13yR2v3w6BCz/QWE9Yv5DctTJ
RSPKzBRSlkml+ligJcgCCkmO2l7FYKZpfHcte9CsaUy+rrtLKj8GFDbSiNna3QXq
zyron8hBdH4VxOjXq8BYB2wArboiK/eX8HTaIN69tF+TZAlSLPpzJ85ey6Q96Zj7
Y5NgwOKxpjejouGuSmigL/d2h7uUtO2eRpO9RSO3f3FH2zVPXZZkOTPNKScRIVBR
wLoQ0ZcCzU4xO7Epopm+wUuc4v2g8CaXmgvlr53+sVUQ6f47wDR+NpGEki6h480m
eAYeRZOo7rrrk8JU/EruWHIvyfqqOAfKlKvxEdVRJJlB31tHcNYC1czK62EWpJdw
U4FB5GlbnNnFEyMSQlBwHNwMzd4/SSTjZ8XWoLlE93WV8UGD7I9WvJMTuFP8bQWU
YTUb3NYYdrmodBynPA/273OoL46KBEhOd+RTfPYmhTB9wRUCoqGcXQBdZ3oqvHik
xlQ5JFcIXrp1pl6WCKvBeF0OGFZ01ZzvFuejSV4BIx8d5mP7ri3JrdmIl3eLf3EP
zPrgrMzi6vkLrKwAjJd6TeZm28lii1vqLz6JA+VV80e1RHAOBaAw1X4QrJkpt+3v
3dYMNnL+jF1vPp6WCIOO78o+xMHIQk8nVc6wnRgZgvgILEQB532fBQc0wrs8qixD
0gb9NawgDMkyyRL0clFU+QP5FyP4dGAHVy2FokVwXArNPqJ/a/9o4rC4aPbbXG8J
EZ2Pgy21MXzBzvqED1nAD/FB0YZA5GHbH8qoGwQCs1Nbv3S4dPtNfYjcab+yl4uw
CNXAPy67yjt7w1LehOPQ6c40UyjUg33wkhUFmXB7XWQVPYgWBdbp5EMhdrLf3dv6
WKmPI0bhImMqqNfOzwTHthd7O1XCWuZZo30eGXx0vIuAiDdR8E4qBn8v/6J7QHbn
Vr+CQ1fumn1Km9hOdSwWyBGM5kjBH826URhNCkUPQv8BdfSND+J8y4WLZus8OVp3
VyhqyyjFfjGluh4d/dxWR+wRzJ94IJlrT9vclH9/CCO5c7WpUEzch8JgvkkbAJl0
45fe08rtcHC7OzEgVip39fNR2yvJVNk0zEHKC4ixa4ie8QHJsFUfCkKtA75yI5pf
syOKcxp6RULOTxaDLSSCMoTkc6z/niPq9Z3+M1qKBLnZr6m74ldO6pYWSu9FeEaM
pEhERN60VOufZW52VUr75VwB3VRe5d44W1aqc6CKIr4zzepAOGaTBxOCczrz0vOX
Cn6LhTl/UQjxBGDUb97vIRbJzRoHAs7CJgDNyZkWVqXNRvmiX27cI6NX0+T9vijQ
a1HqgFmIqZYt/ANMkrs8nNefQxL4qwOoJZSTg02rOe6vLCCJrNESE4JnbnGwGtEZ
vDjU9OXokwiQSyJn+K208HaEb/fkPDWmGN2PVkWSmQhfox/avthLdnTlfjZ3PNgW
arO2BgfHVKhh8ZtNn6hddPQmHrtvyHc0648FSrvsx5scruB860UN+LAw6T/ioPVj
11us90S2FDFSLN4gO0/9VShIMfsSnTiadNEDLL4DuMgVe94m00lThkZTamxI6zWe
TuvpX11+v4Dfhv1n1Y4Bqysnd9oL/PwR0IpmxvgzNyDa0Z0ugUjMh8KnsO1Ef4eQ
d1LXiVFao/mxB7F34T5FhzzBK5cwjvjlnuNxcQrx88FMbvdRBnzC43dn2vN0NpSo
kevGUTYo18np+dltzbpIPyEZJrC/fbR8o9F5I1J5r6ws2XTyC0bDlNnU/1WQNquC
6ZMMMFHPnob3VxIahY4rTBaXsuXhJ2oj9tzF9FKm/9Yiuub3/6SnUTfafhYkc5mK
u3JRlivK2vKioRcWKXpKy6ORdCbKjfpJoffPEHOlAnL/SQWUd0qGDkn3LyLFtRJv
dpx/AZPolisny24G8ytmAxH/YyoBPOiiNKriAospgdOYJHwD7MrW1Wxl+V14i8x1
x5qIGxsGWaSRIA8KMxV+acyuET7UErd3+SzpLkEtBhSPi8dZCzn/y4VBZCgx4ufX
wUo++Fw351JzfYw4qAEm0CmM0Siky8Yy18gGLukdR4X7DS7RXZwQMhyyoatjlRKj
pIZJ1X5wSV2uDpc79niKEUBW48TmyJ3D7pEMV3k/4jptY5ImTRv1tlNfUxl+vuLD
IY3Nd6/HipsTs3ppqiRewGmDE/iWfLgSVG17clrR4HquDTgjHCqni7hhNXDMlEsG
PZZTNgzqA4cxPHm0l7wblNiACW2YMhPZ80BlshwEjWiTyJwglIDjEcjIkjZZwhZH
G95iPoePxXrs7GDJybmZm7wY6GoIslrYtCkfXljPh5XWDfFD3vgutfz3kiXXtqU1
+E4MhYsuYIlyuwDoWjvQSp/TyKKY4VP33EAIsu0TO5geoPeKQQsgw2aIm37Bo0J2
yaML2Xn/1C04m7bbls8RNUnVGXCfDfwJtj4UlpNLSWMqEh1nqX6ng5l0r64XprxQ
QMBjKlxQLU1c9BlIFcqHzxNtcuJdC+N3BJOcbSl9WiGaNa5n168T2KCN1978BoRo
WOF7dSmSiuNt5CQMRjHo7OChS/Ai0h+EmlfzLTZ8JhjAlKmvplpG0tZ8kkyTV6wa
S7wUPng3ig7ssjiTx6Vv4pMl91TsPuTV6LDPzKKMJ9MGXivLIwwlYxx0lny2MZNd
TYRTWLUPV4+46GoGBXFmXtZlwxtv1m77U2IpxR/OmXz+8PrIkNUlZd4BXvGIzyo8
GF2Yz1dcBv1FXe0ahI90p0GLZud3pJWZc6EMriXjgrq0XligpBYFuEdXU0ht0vXc
2i9YSSyl9OkBLYxyB+ZNRz+ELtIB1CgLcxUHr9GDVexROlVylv8lRtyfqqj/mgWX
yP2IMITyzl7koupLw23aHN6UtWjgwLTTKubuUBhcUgHAE+3u0eBNDd0WZMvE0ScC
ZzxO1NMFa3y/bJU46JLjgTsCF2uK9D+thW36VYEsqjVzAamF9N9Mn/FnMyY/Lj7O
EfcajpPFwrmGYkKeWMAeLMO7AlMk9DvY0s7mRToul/Apf4IXhdhMJ8QJa8tEEHGf
z1nqNzprpLIFR77IsNLm7sdowtE3cbRNs5BnOchvRORV0u0H66gG7bX+qO/DC0Md
JrDw1OQMvFPIT9/KEH6vFjpXU0orqttvKu44a4GIT1pRSMXXLWd99wD64xK5blA2
WSd+iyVHvr7K5FmLktohv7xtGM01izx8Jg7Z8FX2ggzJs2GtvxpuQSUi75Ni5Tmn
BV6FFz4aDlpiVH/djw9BHz/xIPjTQdGzW8xhIaYhMqJWAEMH33F2sMQn4IGPGjbB
5T+qzIvRC3rPNNx4cQ+KDl//Un+RwSRdM18Qniuvol0O5lgRdqT+LRaOdg8pRDdT
G4qq7HyesV6HT9izIM8ZNVymkZqe+b1C88chQY0C+I4vWqMHIRDoIcX3XuK7hGs+
k6F4yoqy1hTwVcarpquNYwGU/Mprv8Nuzi91xMBLCz4xHVmrf0XgLfdH/Ek7WDRa
4dJ6ik/m31adbtcxLowiEz8DaxJb9P44/AaGSKYPJerXCSUx1Jbt4CQwfyFfOVGL
nhc0k+XTHZRB74xbR0YiocQf17mMYfqUVLAlIaLrq3x32RDaSIgxfOPKT2cTjXAk
Wyswi3qgjtV0U/IndzMOx5sg+SIh9XT5w+q6P00ii8P3GxgT/NKxSYv9tfS79h62
9b5J/3ja/+t6YpeVBcZ8PsM/Hu/9t8UqO7o9hLRcuzPVA5p/stvqrAsvNE89XsB2
t1caBMmg/h0MGl6NQSl/hHI9O4G+GZSMJcBKDIaZPksFvu2raz02cJSiCmBhyfZI
KBkD/6ab/4Tj0INrN+/28B/T3yg4wAdhpM7B/XbJ4d71EXgdcry+9b19XWegWCHV
ijnBOGfCvyiUL1r2FW1M8A1Hs1n7655Rr/22tFwUiGsXtCF4OIIgkbUNgAapjUmP
HyeFmyb9lrHXqJbD3XM2ma7b7VVigxv5h4vXUrW7L3MBVASH2zzvYW2o4QJbSwBV
1FNMtAmvJIXpuHxFOfk9XolcEAjSUNAHz6TK4a6qivitVLJmCXtr2d6FqvVK7mzS
CayAYw4lnG1vZ8YjKapgO1Uj2B7QWJ0fsHDiKWwVUQojP/7nCUPiEEV4KTZcygnf
BU9UgbC0VVE7XNOBWPjJXVa0Uqc1esjwS8XAmq+uZ54HGS+QDqIk6gSUSwZJQjfp
as3jsl/rvMi//gnF7O5ZgRi1Wqq5y0qT125nQv/qPbTi0DoL8HMNXXZ9p5FaEyRe
tRxETnTiPubozpGMgzDECm97kY3EwXiJAW7CzGCTtN/Kja6epyorxOw8Z/h/O71I
86LftJ0MNkYAFT3hqkHwguhj8GIL4v+EqVWPeJG3T2XBgs2YIOi8d9UZUMcFwYcx
oks+at0bsHLTnzOa4dvqYBtsYoQq5aLig38yI/4EPYaobAD9CBpfUN69Ftiryfy0
qlWrHP5q9e+u3sx4SuHBRQnbozpz3Z9tisHS5FTc1MVX9sfNCC7mDl9nRxzErmDw
Mp3j08BbeBi3SVqduFQDSDyX0P0ZZbrrRtql0Y11C4npGHPc4JpcYvNKzLS+sCDK
UWYkfs8kzPC11elG3gHQRYJWn4CowDK94pwji0knLgA+pvAcq+dmzrRuaj0MaFDd
vUCrBA9Mi1mZLprWJea/DtGzHAGSu8i6qQx8/CI7eo1c30A16sVeVr9XAH9wbyVz
3kPTJPdC4npzZVanV3/76ewrkl9wowd//FX6WjWb98l+WGIIW7b5HL7J5q2WnvyC
Bkp8bXCaNlrGd6ZbvjfQBXMrnt9UjMDrvFBNJOi0GsYLVA4CcCXM7s8AJ75OFyGD
d0JsxR72JENdeLivk8qaDQxfWlbURJsP0Sk4ycV1yOggGNpALIqkkeLbPtOqDg1r
PYp0njm3fSvEcp+VCBq6L3ra3ldmA3WybYThNvZhmoar5LKkp1sXiBHYJvfvYls7
1CoCIHQjCYMX9oJJchm4uDEfmcmbF7iptMoKhXR4D0pqNFa+itW2nehrxcYUnWpp
dXaz8y4cpF3vLY3yPOF4U+ZESFgFCv32/tAwqW4dH1HWuhd8AFpQI60nzjfIYMO7
oN9oIt5IygAFgpIiE7RF2ERLpAAtYf/VAz2QEkTaV1YDUVdPzeMLg+Akfme15ByJ
m3/snrcnjtbmoEjH0jJ/ZyLn4WvH5P4lZwzf3OgUKMEGoVjKFzFbAObIIAkkXvid
XYTKCDY0osLaZ6pDbp5IOt690Dkjb38wY374gtbjyD4a1AyI5cPR3wnVlmIO/Ttv
Q6u6DFCCmDqjmqIAMnlyB2OZZxTiUj8WObKd9v93ztHdbKxNzDYBRRHS5CQXcmLH
yHaIVaY5A6Ap/5+JCTzFKbAZrHf9zELh7wXEmwJuRAgcJjP99/fZUxHlfzXUzTA8
OM0z8Ayr5y1pSBFTWgODE6uuMgINHUAiHfhmDxZaAFDk1C3etIXlaN5r2zClsvTq
ibdvDK81XY2BKi1FkfENZ4J5LyXmXZcvyF49apoZBKlhK/MhwWMeOCkXlJkYlh/e
z623AZeKQ0gf5FgU7gcIuCTREMJbnnCrCnxPXS1APi46rX2LmvBtvR/Im6gc1qkK
DxttiC3gVn5yQ4HWGber59aPHrnCzENdqUHk9K9JCC+gF6CQ7AtNj27OltlIBDBH
CFbPkLlwBZXtqpv80drGKLxQ6mgrwKYArdR4NYC1yuVjNE8YxByBjEhtE5e6tjP9
oSTQ2AXmA5Rfdf4AJ6FIAOBVqTlArd/Tbnm/eTcOXZWEmYmsVbiY754nANEVHi5F
KBAVlSK5eAjC+ignFKsQDoJmtVK1xmKxe/lhHABEbyM0vQW5wwtYibaTYazcFuQo
InJRAT5kXAAxAWuTEyAHqciIgGLKO6/N9WGjDuhFvYA+4cmNt/uRwgYdvFch+koR
FhjWI1kFPSC6d39ZnnIFR12fFCkYJEaDfJrSwzbt+7CuvVGiNsDLV9z9z0jQGT5e
6AIVa3kd8IIAVdD9BwOIldlLWHXAMPCbcXWIHstVdvaVSaZ46Tar+19gnBKPAkl3
B3L6YrEPqIkbTJ/06buwTNTKCMheddbq2pKxqcNvnPGyoiBxEZRUYEWYFYacbfO7
tPP6B/xzi6+ooYPSbijFnUOg5dr10Zjqrzg/A2KyGCJuRorS4iYAsr7Pct0gB+Ti
j8+ZHD56WgRBvEGjD2RuitmBO36BFnLXP0vBpLLWeXp6UsuXX1vG68q31lb0h/CZ
ws2iQswGl7C8iBbyZ3+fU18K4Pd7xF+HZW4tp8xcka/3EdnHxrAMOT7OdMgcM+MR
ETNyDWScbIko3VSzWs8eCG73F3FuePjZZRHHt7Nmk3ew0t4e/2CqVOyZ/vs0uHMK
nJs69q2zTOXLxbXaNavi+7WvpkAIyM37Ue25+ETs9WW3GfhwG/6pEepRU6rzSSSV
TvXiN1eBjdrgdTbqyhnDRdiBSgc9ThnV6renBwfL9FBVIkXWh5lmWVBjgVW8E5HF
jMY7OW/ALBqfpExmku03jxb3mHCDfG1utO9fxx1oUyDJEYQ/Vb+TlTwMU+1nR34V
ZeYFr8unBqZSIN32QHmCAMLVHOPXShZSGZfhFT0DkLIUKQG23dW6uEj0ZpA1T0jX
s/ifCLAsTqCcUqJDilLx3hg8FriEm6sa8YXDiXSgeQS+l9STjm7qClV1vpLvJMfm
/gsq43K4UG+uy22jNbrXg5IULzwL2efDGejvvrBNcyjK67pbBgUJTEix9fQsSyGi
opsMDV7A1/5eDbZz4qPJB6Vptqld3ZQXmb0gv2e4dtOIk4PDYYSIOfeiJi5fM7Nm
KOVmXmMePQ1zKuKXkMB+GoNkB1TjvjcwS31R0xns7qHrCFc5qIFnCFC2xtrvSSao
kXhOLgSX22I5YF58wGhmvVDvVv3kMKEW+wPaAnTR+Zf68WJvHGu8B/YN+qtaCVS5
ASPVbqfp3RgsfnBatChcdOO5bOXeXSovrzVcPlpkW3e4Jy0t8mvKJ8injStjhNDS
3c6gtOkfH54dNNoXXZaudqaB6kYT0HCDVmibyCk/jBsXmYQkWqbHpvjWv9pnsFEB
sZfBhKxKaKDrXfUNzXbieLmaTNBKKnx/tHMZcO4YmUf5tP0vlbdidO502BjZSRb2
ERJqDaK6L5Gm9agjLSQxUCR4AXiDhsfeYSHWMwlP/02Z0QQoccqCBEdhtDZWLpY2
ts9J8dssrDS7/7xdmtBCwQVToSD3klxGD7BhAaLim0kNYqnSkwvH1lniO8sZ2O0w
FQwxAbH47va8/1MHk9XFhcc+PusG4dQmr4JcbMb4qb9oqL/v12ttDkxpnMTiP/OR
E8hmhS0+6GVGCQEvCKXz+zgrMmqH98lEDGpDIM0rTdPAXEDjbVU34tjtxPYYcLSa
j0Znu3uEhDBRJ4tKwwNA5FCufE3pwWKx7NdzDECIzt67MXvU3loXVSTLyZ5mfi9g
ZyQXw2OwwsH19FAUtu+7n10Eq8gp/l77ygpEx6KYisZpH7GPBwc4EO32H9QbwcMj
2jvs4vG4S4plxDYwANX8D2zA2iIJOvW4kuLW2uUFRcWvET02wU8Wis1SIHOldgtd
zBXcxTGqa1a3pZldrWGKgWuMK7b1QKSp2SNnaCfzNKDQl0z+EbYMsirXz/w/eEjA
dX8BfK45O5vuMmyX1NhOeipCt1GJPD3Rkb+SuOBsmMGGNETM6TI7h+JnRcCYUHKy
hzbm0De8PwpuYFpGepPZkWvdSDy0tUdGvHmDZZkh4eAlNLTeu1JCbRg8ngWxbtA0
SyjqNm091FBUyjo9tXAgIrBhUrqeuyhWuA5nP+kB0E42SbWWZATAj9W3h8ZD1YxX
QJB+CsGybnU7cCjj6v3D/kmC/vbZuQdzkJNX0RZOIaYAu2Vdxde+2briF4uYM/6e
ECuU0BK/1eWV96fLL/3EMsYSZ7w43Cy6/PkrmWCkUD+cMkcHuK7QP3SBb3w1Btpt
bFJQK75IDG0AtSkKBB3odeTQgzB5A4V6LUv3lq4JJXuueIHhgeFhyai1q6pmCYSp
S/QGJXC+CxJVo3nqb1iq+BbWYbu+g39062gM5yEoBLxW5w1QBnFH044iTpVbZ3SQ
TNN9mz4jD9SyIRRJsNh3ND98CiaEVHPQ5ObM10NeajguJXs142muFmcOkEMOXPr0
g0ihUS+xAtcazapujyg8glGZeZ1vX6FxFBcj8CUzNoPlSeWwrn3zn/5qTBxdtim8
hBYQFUeTlAIOetdNc5ufLD7QXvoSFk7farf/+SLoh7zxBHY6Q9ZAV/53Y5wtDMOc
Xo/fwq+RKcTLqAAHAqi48XA5cHwyqzyfgl9oiXtd5CIpnd4M5C+9GdBmxt3uhKHu
oJHdZHtXD2nQ4JqEC8YXcTYzTkujWfemFLSPndsyxPYxaa3eip3cE3oKFu/niZuz
l1HGvtVIR4H1OQWBAJfJTssBNaxNMuNvEEi5bN76XijhL1upYtQ50b4m6KA5lXxy
NC8kv+tdaucJ7nLzXhahEnT5RoNQ0l2l7S9QDHQYc8zTNGBNedkhhd3JnTOp6jXm
9I3ev9QRw8kCaBnyE7TY11059Qe3Lunp4isdwVSU+EpFXjqBzvjNnlF7AkPZH1+q
tTZ/xI1wakP8LTpbByugfhi5Q+wVAO9sT6Oubk8ptcorw4HsAAOlPsVaRe14fqZr
V7nbpLZ5eiS62szXaRQjWWld2W/MIE1teq9TlXUMsMpSok9GsQKusc6any5LFJ8K
QJZa7qimeooBf1Gb7SHmT4NipNqbnRaOobBJNq82I1w+up8a/9lp6q7kbNTTinOd
0OzOeg2dP6sPAF+eY7t4OaMW344kKYnG4L4doMqgayZh/haDpc2g1nTI8+Jfj43e
tngNEgb5ks7j2RYbd+/ckPem4Y4UQkLubOaU0fhncfnzOd6fIS0PxFSadFMVuvJK
WhN7DSxsbo2DD0QfYPMUZlCEr38o/MzH7eUDdE94M2UStrbTA5SMLcO77QJGpIy0
u4TS6ic2D6SbN52tweHvr5SO/plsMKiN7fZvEcdKjaSprRGpSItZcTOv124FIfRX
pvCSbWmwFe664ICkHR2lpY0NA4FY2OvFBi6gvmZQRs5ESFMKEhhRZMRXehk33wdP
S83ck9Ub6geccaFvWsGoXX2nzzg5rpeSEPuMbQ7Y324fTDtcWJvPFRu5RrmDzLnm
xNpIB/hK2K15k4EzSrQbN0WB+pa5GUyk9WE/3vQYyHR98sTCv7muru9d3/CIJTh0
tDguLqt9b54VbRKm8xqOer3/+mffJ2uakPVGHwI+UG/1LYrmaiD/hye/FtUMOqNv
RdLMkjq5EMGxhXZFbTs6AiF6LZJkaxraM1aqPjQPpvVcdRXb0s1Kem0rPyQaIlf9
IeyB84ymDospQTw4HfEQVSQq43oPXDZM2HnRjmAiV1qn0+pqO3KPozQwku2FQs84
pT0YKYtcr8afqUSyjeqNfurcKVwSFTcyFlq1kPlzK997S2d7eSSxrCnKvbdz1QBW
qCGDTpDWNvOUtTi01x4PDHEs5CM5e0H+3Jm4oR9kqp4cK+Z8CkkT5kO1Vq8b+299
8+ptBnXW56DH0srJDnJAYUT/8yvbnK8EDIRN0raPijWUtAag+5pEW5rBy0kiZV+7
m8kqMqND2KYVUI6Jw2WQsxKpH+BfPqL8dQrGkuhAEs6nDkqbtZb52nexeNMc3u1z
HONDD6fixcYwReRqJrTvvKjkMgFIYw1J3G2DoDvs/XsFBLU4+/doHyWb8AXmlr7K
PJd2+5rCnx2NE/gKqOiGVcu7goKT1rXBDoHq9q2awlabtzZMWQ1kaai/qQ9+RNrK
BULEzbOeGeAYCvFwhjfZ2urXwyrVoAzKcEyR0xFvSzqpDK0/LPmTjN1LtlN5BVJZ
8rF5omAYDU0qFr5Gk1jj/ruyoGYa2KY3q+ZK5/L9c5vza/ASnU6FV6ZDLz2iKTn0
UK0aye6Ao0QLjnystYIpxwDR4De2UNm7E+c245N2vc6D+HTxdXGbNQ/07TF7PfkM
YNv1wEfcFnW6kUymtH+upzVuX4DRgOVcPyTePc1NCxnhc7kNuUt7ZzddpFws3O+y
xhFL/YEJQTYrDHCPg/5g+Jw43oWGhGNQXEb686hZPBJGp+qYVFY1Tho1MZdhJ3AV
JCrRkmJxW62Xk1o6Xim7ALfEGgIvlTFsvwD0dg0zNWNxkjQVOw37eDNkbAuun8fy
7FLOunXzgljstJUYJDwFtUIyTENQej/BUANdT/u26IKosqxZmZyknO26K3/xJXNu
fiAD1RV3XE+O2LVVsPRGTWhiDkHqO2+gXWRD93o1N46abAuPSZoWjENU9GE+j1oO
U3zODSsmo20hYe4oEZG0aaJ7J7iRL2lHCQKxAfu0IMJMKlX9p3tc1rKBfYJ9j06M
PVMU4mpxEBh3ZmrYDK2Ldb0GfscmZh1LWfMuEhuWwaPebWOG9U9+LfC4XldZ2JY/
l9miIrY83sbb2bRSgZc5oUTDFWrx599qNPu/UNW+p7x5lh/HiA3o5o3WxbOaI6uC
vcDUrkD+uGI13mfliZZUnLOFWMY8l4CqriuskROx2B4lsfrg2Ez4sSuW1BDyHZeX
7e3SiDl4mnH9mtu6vTcKZBYXJIwl2e0Q2BQH4bVxpQfUCYVWMVdplIU71EZvzTBT
GIuXP+9Rw666D9eW7i2JycrAFY8Xjwe1AnAMJTCVmi0nIU9lFiRdwVcB42IJvBpK
w+qjXgt2+ydyccD+MxZPezRzPCvDiCQn1jG/iCDD1P81BXIIVS8fVL+mim+rcWlQ
8YcR3uK0fNm/VhE0dn2Vwh4heFxvJRTzp7GJzvrtLpK/2GEv+h0f7APadPzdulgm
5cVOPgAnkdlCbHjcdUK5WAr5HE8jcYSfmJpbgCnl4RKqBAWX5xao99Z7l7HR422u
zLgIMUuHscmqRezzJIwKPX1YrAsABCU6HGxcesGULYmNO7oWO1CTRLIt5p7GirGe
O4/CW7+ytrve+Og1DNDoFGKuPhAqfy+CaqlfQ0dYZwpMKbZuRWrzuRWhUlWXOjE4
uOQ+wPOL1kWzGQ5RRieKhOwoAs2SiiImiaUUy7bXesTEE+eFNXTHGAuNTvHllm3x
q635G8MnsDLEoeQG1oXSAGswdmkhivpOPmGXiwYqq0NDlz+GKPLySgjc158YgzDY
w9ixvPhHB+k1HC75nLX53LpzCfs3JGOPCm2+NcNkMs5Xb4dbUilPuLykDBltcJiA
nsBMrcTkwzgfEjnqAGg97tyIBS+m8uqJrdogMTRMsBD7FAuVMe3cDcNeu6voSwUT
f93dFsK78AyKzpszeOintqS3VFGGppVjOGXFvrefsJ9uCHtTt5S1kTneO3hndNzk
d4jDcXYd2DzI5NHkhXQ7M8cMxEUOH31TaqmmR0gmRIvbj7usHqIZLZOHtlpAxuKh
/kfM34tkmV7nKLriqHMa/k053zQf/V56HpsnK4Zi72zaKChwagGt5oUMvBAMauZl
9ESsedXb1XcbgaCqPL4h4bIgeDjQUK/TfsKhFbuc9d44qAqTN99I50jRJ9zXckgm
GbV9txRAgZxlk0+3JsebB/O0cAzK/6IfYqGdr6DCtspoqYEQHzb/3niOdOZPB7un
9oAg+Gx+KYB9kiUbBqnN7TfgLGeSyc3/pEJjYaK53euRV4aoi2XGxfNczzQHVHq4
tDG2TOrmWZsvQ2W6+KjiB53vb59AwpYg8gUzQq6J1YMC75AkPzSFmTDEZ8YQG5wW
QWVJx7Q+Y3NH3YNZ4aAwBPJ8ZbWMu7Oo1r5njt9W1tliPvBJCPuTGnljsPH/3vQz
DVy1j9yB8MhTzl2c1BWBdisSaw2PlA4D6b3mJUvfN20nW4aMXbB4qbyLumDcxrNm
ZOXUx95sZXDcNIyUT3KTtJgNV7LnDaBgEEwQB7FNua3KVtBx0ydDe7X97UbTaD4S
0W8jKHKDcTrwsJp0dZDhP1bfHF7Ja8GCkkHrk+iDc+c6pbJ2UVFaYiOLaKC/dg+H
V5L54Y5kCOGQh2RQw9i8ez0FKtE02npMJNvWQ5sf0AQGihQdNzmrM1CWwiMN7oDr
Jg37M/M4JdxTtOjnArgFfNxJL9WaeEu6h6Ll25AGf6Tlr1Ver8JVIWHY7bdfHtmP
xRvWuZtWdyuDugqE44sSi+O8Sa1IPZQny5d0RGy5+Fa3H0+5hNoXCQ2Sh5gmrBdp
vj+yqxACCc7fEquVFwx7eDjRFwIe4dHH2rhB7kzOuFb1BssGoW5dJzUugVM+/ypT
2lYK/c61eLjgKxPjAjaoTWxU8P6XqSY7OB8ho6rLtLRFg74EeYlMY/DUlLWF5e54
9xkKfloNClpyCmNCBH2NfY2fuR/nBLTOjpKpMvPr2kUvGz4/b8tM+eVbcuTJOj7i
GFmY1FVxlwWyA8H6jv5PJexS/pmg4ByNomyIJMPenKe9F+EvVGZlUoqsx5ErqF6N
AD6Lvp/mwiSpDOBIm3phv0MDkdqLvxO9ohsHNncrNNrm+5BLqj9sg4GN4ndY+VSp
q1D26SBAQlzuJGiaG+63a4p72/0MkfOjqchoypHPu5Jg/G3NRlyKUCi0FPQCYeYF
fJcHXZ0QGNO3D5winIHSJZswYip96MEsocyWj4+ZGgaKGSy0yuswjVpYZiyovlzF
89ugmr8p15XyIQmwGE52X2ZitMibwg89ZTsETdfUQCCexiy++U0YFmDVUivUgUij
lWwgmQxL3ZQIc+AJLelTto7FFNlIskSjLJ82phQw3qgm+OdgmuI+Y2daXqsogHkP
o3btqV9+XDgx89C9I54wKa7iLep7VYAo6QKHW192FuCn3/od34GGVAarj344PEgc
5gGYeugCgJqpjgTHz/SuI17nqcJFpxy6Weab1n2GyuRgsh2rQPp/XtYj7lV0B9Bx
/+mmIQF2PxY6HeJrzXrocKhC4UJCDz7rlzouT1AWPiUsYOQv5+RfWOJEPi/hkN6L
CeiEaKzR68B95xLHsFntYaxkDusV0ihpwOC1dBROcMQ0jy+S0oWxKZ873bc+OEFK
5JcmbeoMzT9Dipo4bmMUryf6qkBEoYCJzBcn1h2fuaMOJaX3XVNWx7Hk6PxhjAmb
/GoNFeAh0b6AFW+Mf6SWe9fTkMHzALeMIK068QFgeUIl1lG7ZfjeTqSRhDxOfb1l
acwLTqnZy5OeO5FDYeE4/iKXJxKw2ALtGGECsM4VdSeTWASmK1xE4/Q+xEwJ3S3H
haXdsrM8whEc8CrTGFYQS2+T4Lt0VNg39F6rK53/VpLgGU5rxwy2x0pI8n1OZdbB
ztYU0MGjtbt8tWus9BgXvfZs8LZQlxdbrglwbEyDEr2JD5cyUJvhgNxLU+VpTwnU
wRB9XgeXGtIY4/CNlBApdXldxQ5rybR2pn6d/yLqFP0ilQqaDYZFVU1osBfv7DuT
caju7dciegc88FjKv3y0VudNmd/sObRiNMlHBHZNIzEdmBAIVMyyhC2mUuDsl/A6
iPTpk2ULf0NwfuqQeirKW/Ewoi961WfqVWKFS8du9K4mNLcsFmkW/LxdwVGWaWQ5
OFoQyetav42X7vtOpi9SNhbfuYSpc837d+s7KCKKBZWWEG/m3Fzy9X5JF4EgJxYN
8MzHx969Yvclg3fvSHgiaCaCi/wWTed3NtyX5RRgt4PQjLNhRnKxioPO/3kk6xJm
ERDvJRrVt8L/5mQx9oM4XY/n/FZCMVGSvzEXHkPz2TvJrg+q9T41SF+JPlor8TnT
I0UH6/r+E9M8YJPDHKsIbLnnWgweUi8psptLbIH5N1iEh2RAOJdyHCIKFlQLvg2O
V3cUVM/2GPP/nIl29NDu/efElLp+iEpmtWRAMvGgrpuSVojdG+nB+qJPUUfgOTLz
M7NXPyiP3ivPfVyiZGjW36+yDKyCIm/ZWfffRRxYQKTBxAKMNJDzigolSlXudHim
5RLCLcpvvGqHTGKscQESzzKFod4xmt9yO10pbX2puH8IH7LgfoI870vBOc9EsE5m
J6TiaRPlNA1x9UoA8EkEla+e71BnHshLDjIMuq8CdRGgPtpAZ3lJy0J9Vy9wZHxY
Rk809YjqmpCpn+BSuyx/HA5BgKHwyh32fB36fvh/zR1PxURPEmcwkB6PPDmo6e/G
Vz7iRgyiKEMKpCGcbt5d2FTscm9NseST+DgZ2sarnP3g9vwxgNaHnavZOaQJ3WlV
ulVNaN+A9liWoUalrDjCVDxOWfPO98rITt0u+acrV88B9FAiw+QKMazQBYsyD1qw
1FYhaLR6nhTyrcLrY9KdYO+rV3JdlcLKVpeL0PEJpl49NNEJoEen/mJ72VaSaP6C
cT4v0kV3Ybauu3YadhkLZ/DzJz382BYrGiPxX2nz1R6C0C+5sLB8M0fVJJlA0Ccd
4vv49Tk+WL8f65c8gZex436sW+2GTHSWp3JpgJ5S7Ao2vFI2r40aLyTWFE4mqkDo
L/O/HmKediAL5/GwN5jfJa348krTCDmtbs4+2hrfe6mGcUXOCGNSjEQXJYqF6gmK
VS/kXQThvEcYQbtU4Lv8v+FTJ5kDXqe/7B3xx39g+WtfqZS1iS/eWOG7X/cDE9OR
4UsVIvgr5p2hFM20ak5CH9SwSP6JGgavhvXJy1ttwHRi9efDFhiQ0MPGL1F920cr
n9mXE78ju3f4oNbfWw2Dd5YvwfVJWfy6afYy1fD617DOq+UGOH1ey1ZcCAsvSA4m
Q6onZxhuciU4jpfB1XRwiPLjxwCvNsnZYgmaV8JZUG7C5Y8r045PSwG6SK07aUQC
T5b2CwY4Oft5MitBvyBRds1CP+bvUTc35EEv3aUnTSZVr7GQ0LWStBORLeTh5oh6
kcIjVKOZF+shiS9mJulF+abQjULb/IK1ULELSuAsqwMPMe0h3SPTbF3zIg9naEHl
Vz2CAMbo2eBFxOB0riqZpwlVP04KQOl4nDNsbts9sgB10L1V6/r5j796CUPM3oaF
IRdR1Q0WbwkOJWxSOrjWh2OA40HXBKKgXdYXgj+dW2iGQZBBhGHtUSz+3z2lYg+v
hEJz6AYouI1Bd5MI2z3VBggNn+nETmovdlOYh7PTlfKxptr86vzlZQJFP49ii7Pe
wAXIHPmelE5DwmfDiix/rt1jbSfoKLZFDVd6xlG7wAJf1DFoO4Osw0C38diXRf3B
Z7ogWYq0eSBdImdZ7QN/aWPQQ23krpa1pmMeSYPjLojNw6PM+VXwMxLvsY2WH8V7
iebtHQhlMMPVZW/HaKc33DOVyoZ+KF5Xt0GY/r4AOe9XLrisFuSUYvvR8jjrN9nm
D4Zdr6iAzzADnhRCMxjP8YjNgx2ncSQxx0Z3iscWyTLb12SwN0h6o03qpOG/icJa
SjbWN+4Rc2wnDz3x3I3nT2Uc95w14q4GPqzUkqZO/MS4JS/wOa7pXpXkgkAj/nP1
o+dBotUmhwi2S8YXH5sIRqhcSo5ejqsKAlZ+echWz5FRUHsrAFPljwud6xJi1C9d
GzM8AtjkcbXqxF8Vk5c5gSVgPOpmEBkwmFhIiU+XmKb/9Zr/sAhTWivK2rQGqPpx
8t/M++nM/R7ohBsFXHxXAg3R+Fjs8ZCQkCTtu3w37kOK/uqhOIBXRO71DKx+6yAB
OFaYN7JtpYsJuxCXuTSJdnPQm7a4DPHaBFCv+vgVwGAXwQ4xAYtYMzvyWvgB+8O1
1jZQJ+uLmig4de1bKK6+zU8eqMGSKffax5B7rWFYHtY/UfheAZzAEjUzAEIzFF+E
UnMaziuvgfWpFMAPNqCHAJYRswCiWCoNJH6/kaOlMPZ0BJ2520Kf0BlimoxxYh6D
zAciX0B4FiKl9sy/TvRmtQUMa4n94qzxqgd+bxJ5zJ49fkzoHOdOuxMaoXqmQR2K
8zVYdsoFYUZP8CFzlK/Jto7pTN0zh/TuXvaUdVtSm3wGsTnK0Dx7ViJH3RiYsJ1h
yydmGJu3d1Gi9cTJnpf30ryVT1V5chWXWZKjE0IIgK3zINkyWyBttg2eOalaP79t
8X6bfCpNT8eChuvu777UnkQ8Uv4HQHSqKjUbXfw/F6ppGYzpVDi9W0z0GnmzGs03
2rZFFTTeUPEmcnH45uESNIY6H8TfCXz+GEVida3679enUyB7O19zHUX1NRHVsOMb
HM6CXBTAJwyr71pICy6prxx/8LURirIpO++xSr/Mmr3mFgYDV3zMls9zEDbQ8UEr
tqfJsnRTYAFpr+85uLv4y9ijUi8FCMgyuuGJbyFfam5knB2S1Mk4EqVi/fZGvKlw
/ZS3qQHHeV6uXxQRA/34JFslkCbpSJHju56bCcLmDjBBvsh7mEbXssW/Kcnv/+iM
K6ZFIo/57SzJasv2ukTgCoZqWC3Dxby/nDdkK8ndmENt4Ro/f52bMBjleWZelaBx
uhYxQCf/8tiepOCVNkdWEmeLrUKgT5+FYRvnN+TqsjEfSd/u5bX5LhRzxiHRgrDX
D5TpDE7nFNq+R02IWrhBP1OCsj0giExlqd1yaa83FU+8mWcR/wQNYP5iQkMX+7iO
BjyBkRcQjNYZxVIKIlYUtzGDdp1tbe98TP7JMKEBKCm9VVxu2EaWKbk91pV5UsU8
+GTIfsjX23kk3PhxohJmSo4JXfFN5lxHrduLuL0VobBC39dEh1xv4SRdudA6WDEv
tnaL/aZx8AyQG0KjMTckJhIsEGkgC7KkaICJAn0zyUc7XrHUmTDE0uTnS8ODSHHL
9Uwqk+d4wju6BDT5zXUwX0nDeuQ858OdHehbH1nxLYv1QrV9sGZk9JxFWrxIAH6Z
f44GIYyo+L4YhEeX0dNaYF51P+Z++qiDnxS4AAXzarfsVntXdkhTRBsDB4aly6cO
MoQMi/Ug0sowac9OtHQmd2IoqOm1ZSz9QywJqjvoZoHyYRivoD9mIAtHhSqrNqtS
Xxa4oqpxm1YjXJIiRxQhMulva40uVnFr06LahlvHSvJvGVlzJvPfl/gcdx2gQj0H
sCjoTKTCJjlYozIo/CZQX/5cxd4gGPjk41K7hnZp8p8SGPzp+30OeyiZecOotfHy
ze9N6ICgxWAcCRYqWUNjYpk+ke81kXhSaM0hHReTqy8+cASDzrOjh3UkIbOeTzM6
73xEbEAJGEr2E2BHzEHTQBkdW+VoeqPHPC12klKsZcJckpTvlfCOm3qXe+0bqASG
AXG6uRun1jgq+tXIATv/Tct2r4GGoTAeF8JpjwrW355PUjBQP/GMSABoZpAVDyYK
YT9hjd+QLIlbAWNNSOsRL78EX0YIomhHp4uFwT/+VJyJ2pMBiknE0WOzlej+ndga
APS8EGNPoZ92RskEoJjH1ZhmxMOu00A4xdPyMo7wG4rtJ4ktV9T+sTqQ9/ZwEITV
2jMFs5webUcXZk+my3WiZPGXQVQGjPAgVDO7y6Tg953gRN8AsYuNSFJKB8Nw7iZF
t7ee4ncTMR2LO+8MooR68AnEspGB9jxYR/uSpRSpsJgwB2gmBa6OlDTv7PKedSTk
+YqQsJQbmA2KZThCCUTX+tGjmTTQjheQxkB0O8xIUd2Xn8zGs87NPWGxpJUZ7SUK
AZRdz5EpSwEFLnY2hFDGUIXL3jOyyLRUsgjrlpALhcFElR3Q5Xwgo+zdTyAPfi3I
0SgfdXqS6hUmJz4ZnuXwh/zBr29A2ZKe6LV4CZHs4YPZerVi6Ce2CklSwAzOePxE
DAa2Ds8AyeMm96Nv4VcVYoxkUQzecnCVRWW7eEqThTmPEGHeYldbo1rsU+f8tAH7
Vt1pCoJC8LrJqYZw2rGP5BQz44UmuO4nz0n9FUJl8F6LZK7aLakJPu2f16wO1erN
ZrtUPa65sr0RIIKMTbPza3/+XAPI/D1p95IxB9RxdBNCkf/qxyebKdb1N2n0D28o
BMr5mHDZlGVpJ5/73DQj1QywkaYoSOkrg+Yab4yf5GrNfZhcLkWK8B5NvGBO/asK
7qC66MaWAAyhWoSFhW9XWficyU/krR66Rewp+0eH2TMgyt89W6ti7xMRo/AFA9sb
LJXz0giEnOYOWQtlb9JI1NP4pN1HLyH5eH57ECyMBfI8ZDyWiRdpmkvDvIL9kilZ
6B0AVnM7j+FTFYbVey+rQHkz8pyc+8WWXXVcKhCdHlh/q5D26JVckBkWiqG6nrf8
jzBGLTLGDmFkRafc+YuhtNJuQn7vLfzZUH8jgTq3Dx9ezxZiXGu5eknPXLRHIK6f
Hj9W61atBeZ+vrdc1MNlAZEqtpZQBVHxhtUtiYYPxqSh1ZN4jMLVs1GDms195dQj
R9yVYS1LzPz+uk5A8IIy6knmuEBkWCmoPWHw6chVLcX6VOH2/CzRCXXEd8PbEtfY
mCKQm/Tk3CGFg6u+q+PoKRROn8hY+3WedEG922ZdTFWZHh2SCqlrYKWlm0rSSEZg
NH5CDPD6aOmdZ4BbgZmEuN97CzGHpYco0mJ0CjwTizypnK1lmkBQ7150yD+dr+28
PkddkPu5vTg9W355uZHehtJmXJKBo+tMP7xiPVYt23fYob36rqrKBipcFR1Gk7KW
7sxzhEihnfBQ21opGsv86DapSe01QwvUBUE2MCu2+QldHsPEEqDVMNz/E6margry
MHZFdFuTYAZumWyAnEAT31e3UIgCER5Id1Ul+SyQOr3IgmlLmaYPemdTXN+xNPGV
M1h22m7ZpBH59j0ITl2rviSof6HJ7xjM88SiBACmoMc6Bx6jSxtZeHn/3c208y+9
J390WkcfKMCnbaq3UwsG8w/SJ2r2Dvcf0QcbtOkhOQ85a9Q+0gKLCBfzZ09VZtpm
CPMHbIxLGoWrdFUcuVU1le2ubwnJI7b/VnarZPsTo76KYYjJsPoKXCwLhdza/xFq
3qhVHwTPVkPso9xu45iKz56/8wlGMJgoLAX2k+xBcfSd6Yc6s1qJ8dClI+Or7IZf
azkGrofesWpXJnCN6Qt1OPKI90YTudXOZeDJ+8HlCiho37Ta1AtMyKTSkJwlzHOn
/oR92O9NYzAKNT5Y+iLaG4RX8waf2kxw1YXu71I8T2slLbBkhwbssbq29POVdh1B
PdJMAfN7DWAdu0WY9oExxZ0t5Wj1vPq3Kg+9z7Kv3hXXhEAr/2Og4XyegP0CLMFU
xdRKHHsZqCjUuiAaAEylhlpZWTEcdw/GuNrsmjPmwLXGihkXgDLb4qqijgkPKn4v
TBFgHY0PXGbqQLe6Q+oa5zpIZsar3YlJJFgxYgt7woMqhjus715IkC7kdrn0ccI+
Dr0ZDErtbSpuAWhHm2m48eOLtK4nBDSloCBIjEVWIO0iIah0edT9kJKcgp5+Nk/R
H/b+3l4uXyQwUZ1P4OX/G12/GJTfe9U5cABJxs8xe42gdOilOXn2Cx3yaR9e7yw9
fNzmDAzNlp2FpvWeE8HX6z3KfEzUlA8jL1T11jsO1kZzNd4vehFsJpvj/gJBB3dF
Qq1aMkdcUF8Sv0DJqZQb7pxIz+xJZglEztjTeg/UxiWu8+cPdvPv+wOdu/g0tcgJ
R6bdQ/PJwgqA0HugubLKEf42a9SndyPpNq0ZmvadV2WcegVd+/vdcMYlII9EOSO0
eczMVYNyzA3vyqrX/H4RsCOo94XN6BUeBfcJdOoq0yzupsSAjjWa06JpVrLVHQJ1
YYDbGNdUk3pLulYHpfnIBINrTyjiUA8IUu3SrRM/eViUdH4Pz0mEoc8xS7ud6N8/
AaXlzLXPs4h3pRy5JS1ood10/girAOvd6yM1pVLzG8Mjlr9eQ7B9ZUvLuFX+eWK9
od1hdUFUZ3ZYw+ZuDmkAYDrQY2Z7MdTRZJFti91585uChHk5io959Jipxae3PoMw
JdWTwragy3rJCcTLKNroeZz7HVa+pftRcQNismw03ib8nVdvaIoFMMp0rCwIIvKh
vKWSv2R71Ud2cjw0IUXsQHgnUEfeOa0Qb3AeIGjreHADN4l2kz8us4YdzjUWhmMx
4/Gvp0FtEWqHM/kxtEwtiA51YdKYZKA5YzxJ6uUjdpM6g0e0xUBZNBb7TJa0CnS5
CxvArFo6t81YofOybc0Ljqhvt0R+uUFVkcFxmEfrodTih/uxytEFGDXTk5CT0qyg
QhAKhn0mpX/o8ihzB3b2m6r4NurT6WLTJDCfWW/IGgNAorMLRt0rzFAqeSlpnMl1
UQ2UUC2tKMlZnJyHHzs2MXfTteRE/noDEHSdlJxsPUVOpJero13vCgb50ubwTpMp
aO0RFB9wGs0OG3ov+qhe89Xxz/mG10NxqviyF1+jrQJNWsa4sjs/0KMvTGVyhwqV
K3X8gfsAZ+xbuEdYimSdNxlBRoCewzTblc7Yz8ngqcOA6Ypoz32AbfuA1okb8ft/
+KBEF5BKrgGqBxE+tCpR6y7rIWszYqrCiqymAA7NznxNKXjqqfny/IXQa7LvTaj+
c1QQ1UeXI0PpDY8r/NndK86zLzW9Ca3p2WHcrDRKSE3qAOEYOgqp+tno0BSXUw0I
rUgjpXTURJtkCohHtREeLxZgbIMSt8RgmY5A5NBWSF7hBns7wyXsPKueI9R6L2sE
8vqu+oS6ciVgvq5IZdU5xa2T1lwgyBukuEdB4Uav5DmSv3woD9DEpBRJPJ0LBE1l
utcXH7lE3ngk/yI/5c9v/OAMPafh/lcCJ1tFBd8kIySlo7YGNoSik1u2UpSu8lPY
/Wl4uHY+eYiio4PIm9/1vGvhzXWHAVwWaLqMjX1iEgtmMe1apPLZNMZH8ZCNtNLy
ALTFiHojuDyONUWU9dLPs9yHCyD1ewZPhfBx0KhcvyyIMZKQ+klmlSln8VayVXgv
JfeQ4NNUQMRMr7fSGR7ezcWTQloG0jHqRPff2OIfofmUH0PQafrjUuK9v1heYiVV
FErcZmWAVp8nwBYECeDg6plOkitGOyDjVq/U03FUFIkUJCKRgy0N69+U4Fixu+ys
o8jco4czTn9j08ZXcReNimES5X1AZCWSOWi3OHV6hVb/vLwu5CQE2VqX89t7zEu6
YujyKp1CSg+8m3qT4DRpq+BTRL6GdvoY61DZ+4g1jjL2VA+ltPBZefv2Nwb37hHf
FUE1nqiCb/1+PX1QaEC4VUC0Y4o5cUWtE59yq3NBo+UhYPPNmm5Pma0a8AZiNbnb
A4JpZ7Q0EI00Zj7cP70fYuYhqvm/FhRSgZ4GdygTvMJqUm8sNjmPhay4GqUudeqG
XOzFQO+TFoLqXWI5049/DC3l2fuawDfA7CIqiDa6E44q/Kz4dMEKqlXEUhkI2wM2
VQy5QRDFB+vYGMgavsuxj8VQupM31P4RwRNJby8uIX6BVs5ZHnKHhFnU392vg+7V
JIvbTe/TPuyqOt3lJ+hWzUN1I9+f3OpBkBCvgkYhYdKL/WdQNMT579lf/vRoQLtT
2fPQGZRIVw9f6tkHEp7y608illB0iEoagKWaPM8Wde4jKkOvv5mE8wERNU7kD2fY
dYJhUlsooXpuxI3eDb4rHZgQy0VPW9QDTb3xzOYjhdCZJsFDItJ1wukmDdKtzqkg
x04NQE+3guByecHjTwX6H6pPFBfLYdrq/8jZiZOzu0Vmc2TFNxTo97/CUcu0YOse
IiZ+Saj/jLMKvfsQfMtl7z9eJEeP7O70iMFssRi58nKGUnQs35tH/cHLZqqqG9PA
UAkDEyFkTPPu2OT6fRZG62sR7VxgaBMi+L3U7mZ3g0Hp2PYLm8xpN3sV/0BVxzIA
9ZMwx6Nxoq1xKi4WdBJdBllFNbjToIRYlb7K4uZ57lnPk9gfpfsGQ7M3LDmrSV58
FqISP0k1deJRk+iw7zIt3Opu5SAD3VO/lLr8TULSi6pNyrzgPSaKO0Vu0WARnRLH
Zs//c8xhsOeFd3gvF23ZELDlqhEZ9QKDBQL/ke6GCCEjOisMybsu1djrY0un5Yyv
1rYZTCugNnql7BQ2VOAkdC39yOaaW3UnW/xDIO+KmssEAl0/Uxn7nKr651laVZQG
lLHre18avPOeurA58v+1lzDuLK6UUzHFqdfzfaI+WIdRBAyxze5mg/WxlsYSn949
lmy7mKbZvasOqnOiqv+p4SkOEmAFV/2KcXCgnLbI+5888YU6qydlJlJFx1OEhXKe
CUlcbouS5kyaB8oYS6ojAz5PROne2ZDCE2JC83wKBJgKuxq7PP/CcOOlNhOH9qMU
BjyQWjyuYjsT445S0vnlwStAnczI83Op1DGUcDpUm+VEcXcuz2siYMqiBBrlOgaj
zyWG+IY2LNw6gGldPUoQnu7HJeoUt6vunqTqyPFQirlguFr3ecem/f0Ec73s6mU0
7LUf6plalIma9RIPhMzEifAShmN9EpjxFVbiodH6DeNL3d8v88EL5nrFROz2OnOw
SLJwf8JE+tPmmqfLbrhUUKgRB2FlNXcNngj68N3jf8MeYACZTe/J6F8BCrC3zKJc
FfMSu7zZBvgytWNWh9rhoFH1YoplVf+YCrF30HuAvkvsJOeQ7uz0v/XxZvRJTi3v
b4AgvzHUyF97sZMxiV841EYrTpSYS2EvDzgOHLLuzi7YcMPGLHOGDnWBN1kXRjxm
uJDmdU2w98xiEgBdeaN4WMUJZJgpdfqmUfdOkGnBw8G8jfc2hYTSrtm9wlaoFHNg
ll93YS0Ug/wAiw9EccPGjBI8UVyEaDS5zIAvW5F8J8X+8W66z7uEjJjwlNwDG7am
XG63JT0jKPZ+y/NkK5fUt9oK5Y4sYpoxXg350RLu4UIhdAO7kqrbhsnupiv3qEv2
WOUXR9eRj/S1skoKbgdUCVtSy63WlI24URfT9d3Zz3rXUcd5R9cfx5EK9KMGYlt/
ry5mol7NoT/OnTQ5t80YD1TI3fF2tfFcqMOLdIBW4d4NVj3tXbTrddk5VVsna3lq
Jz7EQtwj4juIMLfk0VbYr50KvbXx2IhytQCnRUdy8zdhdPTj7MT/B5AYqowd7czj
pKhm6WKd3adF6Ti1tEgRsOseqDrMFo5qXu23JDQapj1tc6ZKZv8LndkuhRdU42sG
IiANDVb43GOxPpr5nyqhIGJLyNhaH/cAnzqtqhBKTYs8NXm8y03HZSpzifQC12cK
pLgWVKOc1U3eIefgknnkY5q/nXq/cEXEhnVi7aO1nqRQSeGjIMBxlmaKcgB6M8k7
aKqUiTnp06hU5pU7iXVCEJKzkjhPt64u2SZM7Vi3XsdejtMHEMnqbckUNyVys+z9
kI6d1L6rCwdNmAMTAX8oFEVY5RnEpglS1mvmBwPS9sBPustxrSv3PJCyvwW5oZgk
lKS9eCtAJp7QnPEKLpVXeXwaKNWsjJkxjo5WMzA/w3knqC/vsFbSM74ZmkyR/f90
3C2o0UvZQ6anfhpkfjkg7XRZZ9jVfp29N2121IYj9nZWEJ+ptu54KMimSNHNFpyp
0ZOSL9JeDkAHUZGXhb0SpBI87YNR4GbBBeoWgxSgyJ6M+Ih3BUE8azI3p3N/u58S
u1OXrrAemzMCv8mP3bDwkJHvQEUqsq/PKDnuhp/SlE+ZRsWviJuK04Lc8rNgCLzP
8gKYNNwHxXUPlPVrlvO2Y1B5ShhhnuQAkgXGhSOto4F1nKqwgRkMEKYgfXl/Kux4
EH9V5hnv3UnySqaDsH6cDPDj5e7Wo6S8DQ9zdCfDBSozt0RqNWDPBea0P88c0UBl
eNiGqE0Tubbw8grFp3Qf4GPJcUpDmxwr6fUa7lwcevldk5CFVEqlVXF5EVdvZgrx
sBV8yh3uwoGS5lz/WnmQZ3THvffzkrWD+jZZfLiCAw+BtG1B2QPmHpbLNr7p8zVs
u2Dno8dZJ9+uR4fuAf51MletRtfCjbEH/smv2p9qquaPJ1RdMpn+WgkgikM9cF5/
Qj/+iYPYZiEj7/QwI6CpH0xKgEFcTHVLjXMlElQ3sEzQtue8fZqjfzFood4q54i4
hepsf0I/joFDusTgRM529tQNlpPIUWx7cVzwVx6t3zGlQbS85dk32HHTD8kIufhV
kPvmQkOAINW0hY7M4taKarzMFI0KRxoV7jx5ITvk4OHlBCDP9e0l1fFBvikaxWdt
bbGETyTpqGPEInfir1HUKmFvBHMF19CaERSlBeMu6Pa0/ZXgJ7JMl3UqStPT7evg
0j3zolXD8TZH4ueb7kTgp8LKO71xc8SpsBI0hItP97wg1/jhPlMvUjzH8+wUHLrs
gOLMDqsjfaE3176gKnzVm+sktvXjJn5Zz8W2vE3R5H0Q+Vicpz21j/ljWlPqHRY9
Ud5O9oE/Px63M2buUUAalzZhsUnLOM/wuNabPkvU2XClwj04tKeWS9Oby0RqIZXi
DYTn9BnrS5jpbiKcziREAwgNG3UhP7ip18381SMg/vJ/k2k4fGEcYQ+AI/cQGDXM
Q77KmQAUNCpw5js7qPtzfGciy0MYjfOSxUp0+uquHuViaZ1e6/BGDGHHW8JgDWrN
TnQWADkdEaX3ZpvWNXOPZkyNQLPCHi1qCJOv5g1hDOG8d1jFPq9J6l6Xzeg2DX9g
3gJre4iNLDylmdqqsKYZqfkgVPdvB2N9DwMjk3/PbZYiwPcSdFNvA+5nyG8W9R6i
IlQVuOqVtXtzlXKNCTQiCiQBzMKIIS39TGKU9qonNnLilAxHsHb/Ko0Mj81Z3o5Y
LcLsl6Prln1OFdG1wWYGoNehjgy1n1lDvRhzap/Lm2V6F7G0ddn6jRhiqTKJIfW4
Xur1y/v+uHCnc46yuXDoQd7ltjdBqJIppvCveLJrzEVH4q45AWvO+9CKMVbhqYKn
5zhpqPNEvv/TmaeBxSo9iXd9AGxEqdNT6EeM3mL3L67aV8MoXTzjIEbelH4pOjAv
q4UUM2a/DTtZlJOb4+XN7KZOz2p3Sk0KZF8HMDl+akkpki2YSh7+IXjcn8qV345f
TlW+rgTBQWA/CSHkZRAicBQW4Lv1mRW+Hj5NRqGStqln6OKVmXv23dK2MUNGYnHT
/gRhcDf+W3im3qQvwmWDdf+lrh5bifp4hEsS+O4oXyuvMeE+RjIiwuqV/i9xm3cr
CxDl8/T+vGmxC4e85ZpkRE2p0AafPIP6fpF5yYNsos2EXW92kmzuuGBieG060xKn
vVQbjGElqFCdjURDWefP8avDod/XictamOaIfTkKQ7dCxjLolu7dBWcF19rsXhtr
Z+j3z9gKOG9wHL1GYCtLV3ZpVJvg3UgueMghTrzjNUwdhWofrOoR7IV3GE62ix/3
/HaJXF1xkl/g0z9JCwyN1J4P7x7gRjh8dkrAMJuAXB++6xAvFy75L61/gNt0hUbY
/+G8NnzNjiaxyTwbfUSTEtnN5hGi6rujS/GJuZ257S93ZhF/qQmYdKdUGcLYPzep
5zRBl8SDWtaT6l7dUStdYC28ZGhQmm1pzBIaSAOusJ0rRbZ1EJI0bAsHiKVSOw1U
KBnQlPHAAXpjyETaiwuTMrcCsKrCmLhN16yS4bulBYe3IvA/0/NKTye1gV4sMEb0
VeJeZ0sGN6vJlYjIp6JgMX4ol0SSKGkqzPFPvspfHcrWobNK7+v/Rnc5RzujXeXR
h24vMq+HJNTsYjiTepzY7pQxJm0T4az+XsdK7aWnE+poKDdy0JE0t3TY7telnQDs
2XW+oExkp9D1fjDPpuqCwWH3A15iEL4F+8vGPdCW1QOmW3DdECIZEPKlSI0S6Uv/
tjvK9bgps1ZScAbiylDIgKkHqIMhsVIoyFO2IXGQZ8OtUhNPhUm7WPsWrrAMMWDj
fijycgQXO+dXsxde7v4VSyPAR9PZUOiJNe0+NAs5bBqztm44YPTXTbF+BotZaCAz
ss7hOajYlQEV+T9miMxVufNvx/f8XKq1iF0fj5uk5bNS0qV+O0iLyF9kFCzQAaY7
1Cnn5GEcxhgSJ9pLRHGP13GBuZuQE3dqNktryrg37hIZlkJov7XN/0jJdIhT7OYu
oMn8YJ7jAQscXwjOptST0kjSEG+jyHWk3ydpDLpp0Tz+nyb6Wm/7xnnAQb2dpHtu
+kYgNFgYupIjquU5zQaSlnMLohwccoxRwSF3UX4UYoFx71RUaONIhY9UfBjR+uG9
Bnj6yj9nIP8dK3FMfVOo8AwX6JR/VReCrkF/SgOBi0iPu0QOPoEaEe96mVONS2rX
MSnNumGBBlVN7OE40ffthlCJw1fURBeqvq2JM7pZkZr5f/uBXNfXh0ahWh/HH5R2
PP72jTQcZhcVZ04V/tyvcMe+r+Hrr0IhhA72VUKNwJmJn7+qcUVzbkzxgx4oGg21
aHIFWfk44Hxw/7k2qWBJU7qgJiCL4U7b3nQg4wlRGH58pzaaLR/nMkxC7HnYPQRP
fw7wYKqKPrkWsfqxuh0QbKkMynafpOXPqs24brgRGs6O5Q5QKDie+2DlvaLMKuhN
m+RG3etUMqfuVz8+AXAcFHJaKPUmB2/Jt4457KT4DjP6B3fr6r4qewQCDa7x3A4k
1/F5rxuDkNgeyNZHf86lUl5etXl2BpURGNjn2m3bXEQNgzrDns4MdxUetU7Xwy1O
tSCZUeqZxHEj5lM/afbdsaSvlWrbMdjdEphcvlRgrTQpv4S6eCvYeZuqo7/1LVqw
yewLqP/ir7JWjdyFsMbfRpR8O6fngBx2JdxkFBv1yyHiTUrsAVgDEhK/metGsu4H
dyo5lheEPeA8f9IR51azjgImy298XYBA9NFH40bdG19u7IWXvmCoGep8tq8sAaT5
ompGSGl4zh9iC+mdeGuhmzbLtUsHk8ABuGWXEOI2IqJz+ziIVEt/oM5d7srL6UrO
IdGAPGqfjbvXpNmUQjPOIe69+8HZ4VQN/hdlzPo96ZgAdpb7lOPAlH+0Cwl870I/
dtD2WvXUkvpTrgZOUSGuRJN1nE4H4PjSaVnAJJPkUwU8pMygJDn1l7gcmkYXYrKo
X/MHODwOKv/P7jHrWD8aW544rRmcUQo0mZDpULLfkt3v0f93qNnfkFV3DtPqxd7S
lEEXkOGTseVdRiIzQTxHRIf0DanD+nrLgmonRu0DUj0Vme+YwQJ3LsFlHHiDUpzj
ML+ABeiBTJhraa96mhDdRGueEGLAaNxfQU5TaP1YGvI58DyUKhdxOin9pVZ8eT0Q
eonPGpurdX92HykqHV7DNEbdONUgIqIsYfdKOgqr+fuLgv823Tr2tYZWW/LCRKV5
OdgdGhzwOWJ/WaelweCbr81AG9AhMh9hGvArk99WAHhiBcgGPgP3RbrasqqELzhV
5xB+IbHslLvN/w5UfZxUNxKxkVHZKhqWtQ0fsyAydNcf/6VJul09PpD7VN/YbFCL
6U2f+ZYqGZvQxKLbi+fZV8bwEJe4UMYL1jIWiqs91qQMEpnJwyUnUMVwm+HMhjZQ
1QmxIpSAuHvS5g7Ao6/fEee4uHPNsrtm788AUaXExVMfQTjjQB/l2ewrUXPe9BFY
8nW5TyIIIqVamO9yzc7X/NLEYYYtTna+Kav3sRm+HRaPE7MJeE892R93sITmxpSn
7NlyPcB9kBLdeTLnHtMIivImpY3/xfMlkIZqtLVqRbdRh2V2lA0pKw92SH+XZVa1
x7FDOgyj4w6di1FSMChkonwJemKBXXmNojaOjR5uexG/KKx76wyUAowxHedHJ8Gr
KybrbMZuPDgZVVNXuQ6dF/LBbqf2GmRHifUCRcT3Sfi20TQ+s7nGFIhGIf6p4AjX
ouFsNusSfwz4fMzmqcRpSQMCvhq5cLF/MiiXMnpbbfCSoiOY6afaLT19N2OIzxuS
zppBLqKVJH9faSfZ3Lg0HN3zw00T19HrbNv0ixQ51KyPZ7x4u9Fh1b2qxK5zAlS0
/1aswK8QLQbZ1MJ4ZTpn64mpULjW516QcaX51ZmjA5HHjrCgVOfILbKDrwjoPluM
In5yW3swGCPOAevZWkXoeoeeRP4zeZl23aQWautOnHmajc+FrVMuurR9BgeJQrww
Hp7B2eM4AHnfWSBMVgE6/Yna+nGfhKq1bjSrDrdyA2aZFMqYWTKQDgAWiiu9zs6y
WRdTl+Y0thsuD9m8/GtTwg9J8p0a7YT5+9k+vKtDqGTnqOYMM3SZKnXngedTjezI
tjavLKywmbGY6CjpWtOYkaz5Z9K+KhWOnvwNPiv8aWpFkd3debcOA7cU3EqC5f87
HRkSbjRiZPkw+WzVlH3zq8Ye5O4E37yIMzoA+jNW7nB9u/FROIuVCT6TaAdZV0cm
+/VTYBGe/ODqpu606C1uW2nmV/C69SeRXTS3TZo5nvjuYWbPsd9uXPYQDK6P9ePg
HPYQkK+PkFAi2fh/RBsx5yuGPVUqXsQNVbIOc3dHMEq5lUUZXctVbaezZ+Ce+7/5
CmDf0uv6H3sXIIz8Eaz8AFwOu1M0vjowdodtNBuS7LpqQixipKVtGNRDENjUps9T
7+WMhi2x1xGYcFQz9gcNDxloCyecdma98KQOWqJkZ4W3WpNgWAfeP2IP32YhDyqL
ZqQP6lb59JhAeurpxlfFddDSa5Auzqx85LC0VF8zde1dHSFbGuwMUA/KHNTS38Ac
lBLZQ8RhuWvoN6/VeM9rfortHMDsNtsCduI2UaTBI5hCRK0VAUjPxvDjVNE795YJ
UmeOWWZu/fQc3hjzvYCv+NHKEk0RSjlqwRglFWOX5XsbO2eQS9Xnyy1Yl5KlIfOD
4b1qImwjNc3DVpTZTyxBO1J6zgIwe1eUzmKk1NZSo1uCN3zsH6iOhRcpNAljxSzP
rCB9P3nFXD5mM5LhNNIlYS67CmGyVwTSRxDX7qurbYKvy56e2RQ6UILQAwq1KeJ9
86lVvUpZOFztDJRJSwSt69YK1HvvFHwVoumpapQljitNHefcdmdeXDGJ3o5wUdNZ
fy2yDzPZ30u0aoy0Oyp2KhAts/WXJemIHjRiavXGxZDdGLgWK2al3La7smi5Glhl
TmPrIzbZRAMbyUmALsetK+C7t+cSOTLdHo8Jt4+eyKuQBvy37yQHGkKEDtVz+gLj
iQE3OlSEcEesxTWpQX6g/8zHnm0iv04gD9A/ibKC1ZMsUMYcahWAWahrb2UBT2us
P3pPsQW0qngCAQfSia1AEPaRNuMpW0PHSBTs5KhsTgsXkPAc9S8QF4zct90sthQ8
b1MEqt0vL1Dx0LXpGUcrK+992FusviTfpKlmNw4kr8u8Yth0McZ1KNtQ610aH8BX
jX1HACRTnCPUbDSNfC6Shl9qBmvGOM5vN6Qt9oHV0iagaaiX3WvhZufHijWuT4P3
zAnJyMETIAFQ96S29tJMJ/RJpkXTqROsbWt13Ss4NSdGnRPNkh6EKi6cbaVovXWZ
n914exYKhqZkeYQy/XhJo00zcBOe85gM2tBo4iigwZ2VLKUVSb0k4bwgI5mdBzVX
2iC8xXDpnuJfLZl2rJ12U2LSsimixp3qLnHOX02NHk+QeogVMGV3MAJ1oCtB4LAp
RncFaGp7naVQFRFHBenotFetlgmqMez4p+vfMkAu2Qk9fpvXCF0lKoMthJgWfgm6
XpMK1TCPoESbS/+8uOOngXlHPYRUcEqsB0zqpZAodw3usO06qGdKooV2wncuOc+D
FEATp63cRJKLCT0+JQAtJzvgUShU6o0djbK43WV4d67lQb3mJW42TCYtJU7jNQAD
tIEwLWIPJOcv+FwkCagd3le3sc1L4YS6DdFpHVluT4N1Qp4QhSBuaCA362BayeUm
dwoG70v4pEWyTisHFFWOpj6JpE2VTOPvS8Mruyrbg1xXZlTGzoUB9Bemh3+21Nhi
p5/Sxelsy8UOwdarOByMwRd0g/3ObflQiI3A7HuuTW9owwotPX9MqkOkGAcRxZrJ
chxGTef7vGGtWRKd4+QhVJsSEpdwukoY22HYjT7E6DWN/nlc6PCxoSnSR1iamiO4
It3V9ZEYL/vRPr3nL7lIs4krOlq5vVKTtV90F4hb6ZZ2vglVVFju8/QOIqxRZuYi
s+ZZjtJd5X2rqKhUZItg4KOQ7+fJpPKdRTQFsGrC+6lIDLI5njSD7NoKy+7namMj
T78m8FOKmRRHE7dzs+CDoLEpHWEk9wcumHs92Y17xs6NgX3cD4/zNBOyQ5Rr4gXo
GVD20eGctvxVvG0uObl3MAPjBJkodVDtJNi3Ccgbbfr7nlcuu5xQJfDRmTHCFDkX
WAJFBPg9cHADLyaTanI37kVDw0vdd25ASZfKJNB1pZYqTbJwhnDgYeKDezoy+Uzb
mfajFTJekm4FyQPvTrUiMvORCpHfMDdolTbzPqSNjC7/fxkxdKiDnuKi7jLhWJnD
KPjM4jR8NfvzwLIoHL//Xai0sjMJNeUhJwqRu8TMT4BP3YL4JSOfr6VYgvhLG+nG
PJtaYD2OYkv3QlZW+kHq12Fg1JuEMuMQzuKb2EMCs3cDrq0bMskoj2MbSr40PBW8
hEM+Y0x92olqN1Wim5tmTVOG190eKPYj4uQnukU1uIcwm2mYEd6r7RN4FXlKkD+O
HWcuwmiWPeCnjjkd7XUsHJlQpQJcGCxDPg93TgxBl4IsU9wdx2/Vr2SHVb+ab4Og
mXa2Zfq7vdnnR4mYvXMubEKQh5Oo+zVO5nRr/ioz1N/s2jPlHq61VA7PMxaodY+8
boTTzhkrtwIU/OEc9wd9rXgaE9fznCngC39/3qmGA4YeSUosNRV2KpNfsxlRB1oK
zq2bbG5BVNQ3KoUEubMkc2Ik8djPnh8sjmzwWk5xBvGxACrCWoZrWWiq4wAfi12G
yYk38uiNGmyDT5eAVkelLwJZMA+QM0sOIbwAzsyzSOrlgbxoK3f6uPUkuWYYWO3f
+Eif9L23BCpr9wo3OKOdp6/abEg6fAAoNEGvHqMSTGvhPjMoCEvY4Vbn0V5yQV3O
xihP/IkqClVjN0s7zNrNj9xODzBcJp0auqOKNJeE/WMMKGdcD4PJf1DWojDtNqSX
kAGjSMi5jgQnl2t60nClhTvXLLRJoRZRx/lqxqdYnr1FazF9BndiP/LBehs+pMZR
gP8SVknq8D4P5zv+4YXvlXNFi7PygOI77mTs4l7dZcpmsd/ZjCWHUMYuTsFXpvVP
rjYjw9ODPbyZGKn2hjctiKl/NTqBwdOlfo+/bxmfIcSt/4V7MKJq+uISpu7/JXjf
xqZl0IRNh1aKWZWbobmQCet9dM8Ritb7SE2XDEjip9f7YELwWGH8LVSGgNRnEs4a
QqiCa3avpwLgfsjWxcP8MGOxPRex/xV+ra+rELYlgQnA+87TlJIeuPYYpXI6hZaO
p7z3VjPy9xq9TB1iY2gJjGeOtrjp5PgwvnE7StX53gQXzzkYfXq5Tn8N5drz7zfG
2ZvC/SsvFfbFoaQc9Y0WWz5DiDHF76zJPgjuG90i2IS4w9Lr0reJMjz4hRuF2n5O
mXi5lFr0fvzTTnmXpgAbFcl2ZtdFh7BhqxdAHfiY/qOL3QgSM+h56iioZuGDwAnP
jvdSeOUUt7Yd+QjyXRYcn94PKkkRKiffVr9WIl6V8NuJaByoY0ZUTsLDRYe9b25p
/iB8mOXbBi+0lsX74235W2bEtQ/4crt1vOAHCdSWBuyfSBUAGcXArTejloURBMAc
hCEdGaFbEN5m6AvfDEWZaI9qXSjsDajN3V+/AmDbMGhulT4cvggNtfAaFOanCI6j
P+SbGuAUJ/TNylgZE8WUYRfgxlyf/cTJOXf9eqUA6n/Pv0YIPbgUvUXuuUuaK9p/
Ae9oo//UY6raO8QcEJpj7p0pjoXYhW+euWsPoxOB7mPUnbvIwfYSqZw6bzflu4hr
s4rtwf1qv7h6pwW3DqRGE9Eu+Q8w80++LDeIFY0FhfjWBmbiaGyiIN0ylijkv3Mg
g54KGHKFQB8/RbWVpktl/3eJ2PGBViqKBoguzDvrEaJrSBVlUVC/0fy0zYae8FHg
EqpMxJR0t+QMSlqFQfdp6/UYZ1tTnW3KeZP+rKaUAjvtgE9MGBYJ/2uS8QE3ElyZ
2aLwkdqiL9BP6bWp7ChO4e/xhyk5b0GkpxrU2avMdo6ew5KzSCVsLjSkO/vA6HGW
2RESQFe25EA5HVCaiOXSDzaGpx0lxFalP2UMddI4o3My0A4xEE8ww7n/RP9NTTqx
TD+HWo0Ae5lwrQgEgngBe8/QjslcZa/CwtW6OYTBNqEZBQh0oRH/gAL0kjftKTxD
A1F3/I+EdffkgmrWnF+M0Q0FzJ7f8hRCLoJua9VFsz8DkwA4sMufB7jP/CzgHNId
FuYdENctSOVDVYk3s4vRBdZkRNUYs3B2HxPOOLoDIV26NoLlB4UHl1UzVgRxCTBL
uFTWzin1Jsor3qeHqfUN2Bpby8KSb8Fn7tejfYY5R6KXa2NXzsCsQhHweO6o1HyO
GA1vefKOPA1izDt1E6bCUfCajTDeGpeAjTAKrvlH4QkJv6KkHOoWVL4G8qP6hyjq
itTMEq3pFkEtB7IUCMtlYSKFFRKS7Yas/4fRUS+x8nmx/SvQcIK4rmmTKf2GsUeZ
v5bTwgUWfIMN06h6xV34HQ9MhOVcXAA30a7bTa2kCKMs4PQiea+BUpqbsJJvII+D
sUB+3foOq0y8kagw58rvGF7ynaDfc/q9b7YLLDFQyquFbCSpRkfTDi8i1RMa2gxo
xAhAgO9zVeEEPGmvvAbG5/N9lDwx3M51jxbRNCRREmIHpOGtmtv2A7vET75Djx9f
i8NMcL7j9S949BskWAh4ETNAqgMbpPgicttbVXuugsOhXspeSL0EHUJc0OLQEeKq
Uq+s/I/gopFFks179+ukigwgFr+sg1ZwcngCvW0hg9xcAQGnAIbjXGpVIy5ssSIp
EUSjafWwke4ybmNsbsumwLLgvRL63CK3aHQGWQBMZJEzMkbrfg+UoLifs0UiKU8B
nvnYRXihqD/kj/8Dh8GaTx2TqH3+Wqpgs1/187qZI1vwQXw06CPT0FWD4uPv5Zvv
FnaLUoWeSm7vDjHK7haMGFZsIL5oca/d2x7PTlO5+j0B6q0+CvXHTxWKXKOjz/7/
pSo9EBLNrElhfXa0oIbbdD2QxXS0GFfyINHWuEKIS2Ev5pFCAbEInbu3WlIB8Jga
hg2X3Tb9fNQWCXH9Wd12udvPAKmfFguQIgVFUkH4m3G/uywmGjdt7US4lPum+mo4
c3LsQWzp4f3xMrwPbssRYNyGQHhxFne4BxgMP2T5DfuudPrh3nNvPRhKexc04oUu
5GgGu80/Z+cDdWN3WsBEG/iZ/T6jaOQFjwf5D5WrTOMgue5tLHSFasaXHbx/fKZv
lnV0JxQxmbs25X+72hWTQs8d1S89Hjv9laSn7PDJmOyCH4gb/j+un7KOmI6WHjnf
TsZDn8YNQsZ6w1O/JkmUVroyMMnpjkL3KGyrUvzaa5kUXP2ZLdEsC4Sfs7Ej/UPE
Aa7lQzEjN64YC7rBSNUXGgSQFSnGnS6MjayIiw7Wg4za8Z+LeDq9MiSC8IU3XEhz
i8/JYpsiIE6JPMTzOBL8JV2GBjCXdz9ruy8whDiE808QbVUyDBDrG6bh+kRHifh2
68jdjWnb6N5PCS68VWQLAEoZqWrsYMWI+lvCKvEGb7m4W1rtCKxiI2DVPv59eTTk
XOYX4UljFs5IaNJ7uTqPQx4XPGEbgzzy4EnZDBOsRmTHhRnElNfyuhhBsC6TyuPD
zRrhHedorVlx6+hkT9IBMKO93R7yVumPc4tuciXqKRtG4Y4AD8nF3GFOJLrY5zX5
aJ4EkhSj12hWYHtk3hsbRYmCaaaPPsfdIjSQO3VFuIJhzWbQf6rrMlsSinOOCrQt
FCUocEbShHGc3hnjZnlUw3RF8/JL4KXpGLNH0jSowNM4BNPTSlvTxMyArkTWCcO4
1nnH/bIY4My67hWNJIUaUQpquDNtKTXMfo/4OatjOTT3Gv3wWAo2H/Y0QmhAACSq
RMQv3Qes4eFMvgXtgEtXG2Hmb5mFh/wdse/tZtIsVz6QoTM3B3Z/FAvy42gvUJ34
xPM8CSIb3bS81yOpoKiQE2P5l4XqdhWIothBybkdb32x3dOPd9QoeWZ//45pFXR7
MEZQV2wEnuwTKLDa8edg/ifH65awQ/WUUnaz2ERHxNdAa5Z5h+IlhDPec2LQAdxe
HWvKQeT5SZIw9H6hwgRCRoKcOqNqOHWLDSDS6wOWqx0Inp1u7DaPGaz/BJMkSLK5
WsQWBuHvCw18mKBWypRaABWGEMK3Mru4bLupZBBEjBu+evkVgGecMsDgAqSQsDUC
wqCTl4hVi5zBKPGeYjAnbeJKsCAxawuSdf8nBQzwWpdfBrgIwSPJPdEOqMK33rq2
USsA7i7oW13rqcXxYLqUogUR4pscXwDd+QOPlaVVNgNM1IHm8qde4frCldgGUZdw
BfClP9cGwO+r9tGjwEF27ttKnFmx+q1u3oKVZNBxZhoS9rqFviEz2Ngz9xTyVQa/
bC2chpLEZZk3nxbGkJigyvc5rq8GVFW8M/s2OB1aMN8s+eDisHLAL9sxBVt1ba5x
VfSEBWjVmZRWc3U2q4hQ1pMB+vwh9nfqhn4kWYab5j+xCB3LCDVL8VHw0HrrzXVn
KGSS1Pv7XkSiBBR9WIaQIm2JPB+QPOUcfv7BTyCqqkWWz+hHySI0UHyPAnLzQz9z
o+A9NkdO5PcT2y5G+gztDehH76k4AGtep6SFopIKzIvHNZDv7cEwM/7qRVlfFWqm
MngHEbvr9vN3Zt6VN7yDwfievL6Lpl1zsgThCdoSe5dWYVXZpAsMSU1flHThCyNd
7rf90Qe5ryJnKwXnJdnQsl6ZezOpWyB/1Iro2i5mrjO8nZzOthpGaQ49WEFd8GbO
BQbF44QezGC7RMOMdDco8bZARATk9bF+Ket5OIx5veN5kkMowmvxII/ChNrHyCAe
RdxNzDXsrOAjgjFCiptURX0fQrO1jIjygUOwrSYH4grXiCBAx1G+FqraP4lB7ggb
y5dnXcCJYedd9C10Zo/T+fHIrwMWdFog+xbNoTTYQ8/jCU0DUUWWDBsxdF2lJK4D
4G/hnDWSufwedl8x2kaD4unIttntS+DLqEGHl0uKcB55ZGlKN2AkLv6f8/QeGsfG
+tm4INNd8BP/kkrlquv0gB0T55OCrwBGx9GPdQh+JtmzGbTqCFmR6GG+wICWyFF1
ysm0z+KE8WIqJh2pzxXISJpvZtNZupA5buGYwc3NokaXG0PFzDD2V6qjiirfXy1E
msEke6R23U3AwsLARajbEF4W8ACzFQHCElgSGPNazhudRwS1FYGyVEGgfyqofnZ6
WFPPdbaYeEGy7NeWCumR5YrBpwWjuXevVmWtRXZeh/c3zejmBoqdUU5vu4TQk/cW
Pyiief4qZAq5hDPKEcQ/vKIHJLZhjT+Z4UT8Ce1A1GyUFLNgBEIPr6K7U9gn/YZ7
fc9sfKJ2IHZmsm+wMh4C6+buyExhDgRtfhw7gfmfv8FHVptLkh7/DaI/9O1Sa67B
Ve8EZRy05s+korjtodXhlbPmehZEg8k5JPdv/OsAzZkqb4fyEk4Gri72TySteklq
dBILi2NSMIzWnd2a1Gjw5ODdfcQEViEvyMtBkoEfx1GG54T3hvPnPb5Zk0M3rGy/
qmgK2QAOQCPddtFSICadC0PY/5fv9fk4A7L/oVlD1WRUDLHTPl+SMovaad8LHWej
0jPcvkDb0/aUgQi7N6qy91V4xNHw08d/1P2zng6gTlNrZvuhG4OIe16e8GyWJvwE
7usFPRzPf73aHVLtPjB3IPxLkFbofjqoXa4TBFQu+mVYtn4fJfyG7UU7eN6o4rWy
1O7N+3qDDPZYJm9BoYo1lWGXpcid8P4i3jymFTazqGRiiSeebgtdzBrD+DnhfX/1
8KBFH1Keztp5xEGg2SzrF/mB96zacikTVicVNFgTeIiQeBCWWMEL1be1/SESRxy3
gOAKU71HSM8lZ5UlsYInN1R+tuZMLrn0OQGyP0P6vLiiD5oT9DMJrStObuGjoNkd
kwgiGiqjR3ysUXVP/u2lVdJUxn4M1Si3H7l7nSL3K/x7tdaYzE/2rswj6nKOJull
q9jbSZ2oG4V6YmceIXiUQ1zVz3mWlOW8VrkKxFmEnrxZ4Ao1lCnJD8oaEWUFoAJv
Y4DmYEkFszuVdvcQn7WNmlxL45gjRS+NLErCQyAKOkVey3fImT4STw1utmQoU7dq
r6XMWnN0iTSzndIALvw/9KbQIvbE+Jiuo5Zw/i2Lrv5x7IKvNaPtRC4VInJA+f9O
e8ZjGlEXFdN6P3RUae3Pr24IqWDBBg5kmgdTwDtbuR3HrLujybSg4cb52jm8BYUE
hcGjITTo/lQOZ7d29x/AAo5aN9p7ZSk5vETumJHg12hoINaxPCrEepOBaDwwVCqg
pvtuqzOA2UbubtNIzoVUR+BE/ABPfASqbUOd/QXcrPGM10Yry/mNWgVQNLyWr2FS
jw6jLtOKzaQeUrkvyK/Qjzog/8EyA5lwUMhoPWTJYsPQo0gTpgRX48hrbbVSLdub
rglrwVP07OnjBdSWtSD9tDxgI+XflrDpE+zXrNK9WEL5YC6F1AcmaoXvyA1JM01a
bEXPkk9sjyj9VIqnm4DFz0V6rUxiyhgP1RrTzqV3A9sFFX82cu9ZgtAvKTDGGuTx
MpXq0K6FgdZX8AUBwloyLSYOrMji14rpv2A2ubg6zNVStVZunkeZL47QzV+URjWX
LIuDYLaIO3+NDzlrg80OwFEII9YEdGgPLdCcwSOaE6kwUSX1hkVgUgUeqqfybRh2
8/bdPQFezX6qC4/S1HtEj4xjZELFFa1RYf9rWHY0cJKPEMKi5/ajrAev8DhiQD6n
IyMdUJUn4xgBZ6Z3gJIHf1tpWCljvyIxKuCQA+K/aa+WdNsxh+nevNpA4VXqwpku
DT8sT3pUad+10SzDfpvouaLjqgEEY0f7sAW1X5AfyFCcSMQm191eEqrmuFHZDQnR
gZ9WCg9j2IMXsS/4ZYtIt11tyek8UlVj5Izr7nX417LjmOmENzejqTPbDFQn8okt
De86YkXG6mITVUj6+SZRe2a0R+D4TfFDgKvUfZR6M6sbamEKQTUbcCE14mBJREFP
uxRP64tI7cDtZKAE/WPQVtB+eq9C1zekwDQMluLHt4L4uaDUQm5pyVN64c6WKS5C
Jh81iNUHVnY84a53X7ZOJ+iUeZ5vlgnmQNrFRtCaytwHii1RF7nsdNzSk4WNnvHO
Ea5itpyXIyubnv2et1iCHn39Fb+XBtmTaJ5BfOOaj/Xb3gP8i+mxSibe4uIITqjk
gQjA6gf5Xnmvb8eDTssI4gAM7y2erseyl1TGm8zd9NRKEOwSYhSVBQZfzdM5sRx9
8pa0k2qvMNT2hF33WVD2Q/yC95LXl075mNZEm7r5K4081Aq7y/J++bZWFEivtb4M
zmjX9eEV96QGFu1g929PAzdO/GGr/HwK0JrCeEoIgwEa6abUMgvN6nJ0W96yZ3HD
kPiWodWuLrlET7PX02R5SXG1VjU/kbcnXtnp/Ap2eXLSutqZT7keUSrLdTUQvMIQ
3Cna9c+3YRI4HJlhicjkLZApBx2Dza2COQjU4ez3xHlHzsCBWjNWAnwgOr+OV3Yq
w05mMxdA1Jvs7KxjBmf1PT7jGfMkG8Gk5wnzBlRmAJip5Yn4DnGCIcjcVlXu4wj/
drEXSW8eYszy0lbnOyN+wY9giBQcVxJPqa2iHmS15/YpUcJmYltO0ZafVuSjkUtH
QyEZ/u4JEslfKWkfYct0Ihc27gDiS3NdE4eied5LTI47q8Eb7ewu6JkkutNFUA2y
HXpfGLVWNzGksfKZ3K5G0/RLQEWIREc1NqKY9kqPPSb6QPLTUMqsSmmz0n05AwL3
z4k6aRDfw++tpEgMbp576WXFPF31fd3+LfhD3zzPUxzN9BUqBUwYfShoyh08fHnR
m6qIQHzv4h6I8ikZHkraYi+uH+I7+dNlps5A/PfpoRKuQdcoUyNEMJgIzbPIEqRn
Y2suhD5PDm7+VbguRJ8gJjt9lUe3LnS16gM1wjn6mcgyfA7Nx+aWgtqYWPjSjiVV
CX6IH3jGpZdUj+mZ5PwZY6zdhi5qvNYfk/B2Tu8HNzVHwQKUDUcdtbnbEMOQnIf0
IYU1c6QZO+8DU8bxmUEp+ljX+Q3v59uF+xkQ8RzJdW7UiNuYi5V1olqbUwEkI+Gm
Bf+YvTiwPQZ/QhMRmryXNERb5+w1SMkJ8KSieAexlW6DI44i/HV4BqS+eH01T/OX
R47PAiNHhtPvXJuivDdcZDdonKaHKD/Mpb01JVpyCWWYg+IjDRjZFu+8UejpZyeQ
68l1YopWZk31xp7TSpMjGsTC/PXpuX/4nEa6lXNxN6XaoccpaerUdYcceUcT9QUK
UsiXzTMBJHrdzjBAC8vYR8a5Ofy3mGHrlMsVr1yGV+WCYzVmCy5Yrg/NMIQrMkYd
Fk13MoZOaVNa6KuMouElQhZqyXQh/yPBJLrN5bc5idM/Y3l/KMjQ5PDrgO4UnWQc
mA3BSUsrxprX1uSap9HZU+S/KqlBEl5s8nEcWl6aRG6l9awxa2BubiRgx/6MOo6z
u8F22oANw2joZIFlTg8LozYTyLaCiJoFaPov8m53VVtoENCoxFp1McB6KFqLLXT8
03KdCQ6QA8zoQ9ast51vcwbCIyBA3vnAf5T5/AiPY3phmpZECsTx1KTlpW8ueEif
2c0AIipM2Ua6gyZlpSxcIPCAFRt6fk4YV5lCGlW/CeWdpDRb94ickVMF3sFawB0U
RRfaI6ZClnOICuUPGblBhYB6J+2IvgPs/8nWjur/RvrptjbbDkbWsPehkcQGpNux
/TcMrlSZqya25VPH7iiNpUYbAAwv+IIpEil30QatL4PBZgLekL1HBKZjAlS9RV2/
Z1Je/+86cc99p+Vn/UsjxaeLH6aQK6w7UL8NwbH80QKAJqSpjczUSqj4ekbu5zeV
PEmkAvOANiqpVgmetsbw83jorEmaVm5ojrIinrn4lBBjjwhC0MFnsuCmnP3IPWkl
DZGqS4Dbec7Db4HlUdJUb9ZDNMW1Byz1L/ioL3dTPAL4zh3jvtlLnU9W4/WY7NHI
G6bWswL19Ep4U8TgnlrDFuz24c0Cma0UM9W1V+aemyxdtx2jMJWD30BKseg4QHAg
zzp1pB1EHizXWkIxYVfl/CLUyacE7viCdtW+67ER65V/uoRIlVFgkSM8CiAtSTI1
azUFMtLaqU/vIp5r1b0r/Caw+N754vHhHFA10bqZyyqqK6q7WF/klozVBGEAcV89
BycQeq19mntjHYd87rX+BzK3o4i55xzkLezooCD4kltB61pKrK3fvp66nnKvt03X
c0ejwYyjEQc1OolMYYU825kwQsbKjsyxOUcJHwO4oas9gp4sTJsYcM6aBsvr1+bU
xJPcXPUGhMptrfG/T9yYyouX9c/b8NBag6atu7A5DSfpcpKYM8Xye1tZd+ZcgjQt
j0822YPkvgdzjaPrmGytgDdLjnPc8Uuu0rRfO1RqHK231MQqkzRSiXhu+ID33/u7
l8H0NjZY1dRC6or4iYp1PUsdcNDqSOa1Lo7IvG2LClF3gAgQI6AHB7c8DHZVktfU
CL43IFHDr91PLbBFHhihXXQqkCZPmHbh+rltAd0T3r5sO6ThPh5VUWaYYxMWDGXm
VuANoxUQMw6YQzHaplYAJBQc7JFc22bq1KuR4MsMUVd8SsY+SaGk/LTvnE2zrUQO
eTYAD4ki/9r+0j7JI97DzDU1TeCefIbiIBOTj8MJhIZ8/nOdt0BQ08EHHv2pZnWX
qg2Q3qFuetUIE4rLKpbxbcfRDR/z9W1XSij+xtaFYfTfY3t7u7Qd9vZE5kjChpTb
2k3kfcchXJT9w9zpQozA93xF0/DxljBx9dPWkdB9tXX0srAIrIb5pAtYZVZS9K+F
4+H3QeUj7+U6VDo4DF5M5efiQkWglerfo5FhChJycL/VL7YtienlQorhwG1+e7QZ
Lc8G14+5NLO35bCfewzGRSnUAOEB4CJc8eBQJaam9B1Q7a0v3Fv+d9dRMjxbHckZ
k3c+fWE+ygV+SEqKZyGTaDPqcMBIzFQFpiF3iEb9N8hxEfe461Qvkfh0CSkhhutr
Ujfky5+JpI3rBIXiDg2P/Oq8OpGRB66Pw2q1RAZdfozI0Hksg7FGIV5v66yVo3Tp
imOavAXpnsx6FhIGxLZ00s0pIE60S6eIK837yHl6CcbTNHyW2P6rtDh3yVjgQnBq
Xr1W8a+ETehziefSX4ZkJLzlWAbQ0YRSB+SkHyoaGiLQCn+cYVqHiexkFZcQJ8AE
uSXjtnF1yw2P60YVvDBZIrKVhiaH411wPDNWaRNcCzDjJG2N9zfJD3Sn0oXnb/yr
V3BQHImEUHurIsZckabUzhy4BkNC0XNkpOGyDVS2uxIAaf1FvM+/iij7IvF70XYM
w5FG3dyANld1j2JIAOpcp8MYI6n1QJPgbpRNeEDgzYhJWZQCZsdlc73mOGU1DyOk
ssr6KBviPUz8/dkN3+0d8RJX1hUJKjLiU9bLj3WYKjxaRAc9PNNDsHZ+t1K6dxwn
dDjVyeRL83sWoaI2vMI8MSSMsmNr7ubBp/JQBdpAFCiW3zRf3LWyJyK4CatUopWI
SbreKTKdXfMM4DW3oC5sx1IapPIWTFs4ivzov6rMIR8PMbnlHL8qi+XcttrAJjjb
5zmk+EfzNU4z0rI05RS3SK0HXYEpks9N5Rm8lorQEQbG5RLvregg/1NqzbF8FVoC
gpaIkCoR1RNmamNm9ADQEpfeIhXQp8Q4gSHUgusBhrlhcAXjyXVL6sNW6QId7IUF
iTl2wLWqNM9PDGkcSiirp8zH1+98FF7lyVEwWyp8u2d7MPMvhelKOnsV+HKFxZW1
z5gQMTWmOg7BBo0ALHIY9dZfoA4z6q9odjTJQ5BZwc4mZSFaT/W/Q99A4KcRJNVC
5gxap9XGd55lnIpyKeC5XThSodmG0g1NLD0Gv+meTPpdeNjXB0qGBNS8t1rPXANg
upY0vzo4GclYZOXFBGidXmvLPEGFCkZ1p0pAVF95AfFo8fLDELjJx/i1/yEmldS4
NGTKcLt0jaaAqcRXCSTAAh9gnSvUckIejmnVl3O/yt8Ydu4ZEVRTewJVK+W7suJ9
utYdMbY9a9NOg47EbOIJ3/9C3x89PqtV90u2CxDqkjulfVu8VM74k/CZ40q9MYlW
QS7ZnHa3tChVuko6lIFSyJCTiHt5QXIoxMcttcWigxilJSaOeTHmhwaQoPPPEbFo
/fN24i5eXo3S5maPDm7LCadVAw9izZOmKLoalbKRc6qdYHsyYoRZYaLg0B8aMBfd
k3knerh4qvQZqTddFMx4Ass6fRAUYoWZvAHb7n3UlSDRa36tRwN+BVM193sRq68u
a4wLrCyCrzYyAFFrmsyfWovtr9wXzS9Ip7FD4+jpK36MGo6Xj7B9F4WSZ3YYKnaK
gdRjNQoFwV4AjcYbyM3bfln10EF08nncNFvYxWJUMeTZiZjOYKGgt87sspMrYIcN
l4Idc6fSlOrofB6LWvbsydBjv02nW/AlJRgy7CsKBpOTXqLDPWpvnZrawHINQLlU
sZfiuSaIcO0IIsFXj1ODJiXs8zM/9gLyo43sO7FoSSuyzQVgn+MkUNgVM50Swasi
N79WL3eESrhY0c5tA54QyXVlDxwolvC4yfpbf9UoBA+Lu3bWox/vhiEj50wF3pq5
uK5s0W3XMedGzTadHezD9R7bHVWfUOQMv5qEi6mQobVBB2lkUOF/iXtD6g68mVbw
rxzd9ZuMKfTf94C0DyxsnF0t3EtiBqaEnsus4lYf+5XoZkk+xtcAxhDL47rLCvU0
meWKSCIpj+OoYa3LZYP1ITAjNCJl8o6Tsk0UAPNP7Z8oXdzH65z5tG5wt2qX8NWa
PiGFmege55BUXf/kailbcLXpO38S5KdKW+QIrSrNJ4Vusu0lDiJr721Pi93h6hug
/j88nEE8DhUTZldmjpNVL8qlC6RFwWkXMz7Phiq/ymVV40/sYUPWrqGGVAIjztC/
FVANxmRHzI53O7slaSHJJcWK3oaeXf6kJp4L4m5g5luf7pCQKnPL7xMR9koqKxHT
ZJrVAtLZurUKqfwVNrB/vvH5FpqMWU27FxNbAR/obVUconlMNbeRR2N7bnMbLvmU
YLbljWVI8mbuLwLUfq3n+BkWqVzvMzEgOVuRu5I/9mhd9my9uh3jAcA8TjKunmk3
whSzna5UIn4kxz9KugaiN6IWJUtlZsxDlu6kqeV3vE4gx6NVsCSpYSV3yjXjyEGA
kEuHIUjYbjcmUl+dZ3pIVzA18bWdDDLf6L4iVu6Y4/DRNCunhpOyF6K2WaD7DPUw
7XpoW6XoM+YetVsm1JHdTvMaE3xXOjAOgATzD273oLCTWh6JY1cT5SOkXTOdYash
aRb7AN7RN5Sxs/59iZsdZflTyzjm9lDi63Qx8/wNeYi/orGX7anqVRu874QP+MTz
LDxsidfFC5URjyGi81uD4ocMnbb82fpiw8n3WeBXYDSKe2DPRf2BS1wu8Mzg0AKH
xw5sLvd2satES6U+mpbHfS3Ej7lClqWbsu3NiPFZlucYddDPUdppRuaiwG7KzlcH
r/sEtrsh3FdIgTUK2/i9zlw/DH16mMyq7w+IETiJ3NyvJGW/2/GXqJ1b+MRfD75h
H5cVJ4A/XjQEWlNuCBSoSXm65GPVF/CqM63WUSX2cDOmzdiOXHNIlCteMKBTwI7u
Z/ogYVQ4ZM2KiZwPNA+6jQXrx4Q+a+zG+r0Y9tmT1IOjGqnMwzp+tDWnuYcOrdqi
oqS6zKa1+zqIX5E78g50UxVT5KojQTTMTLqqW7K1uGpltI2wvwrHYOs2QT14WSup
13G4nutrgO+lzxF2s+qMFbfw7MaYs1O8ceINEiKsvlIP2pI9qlWgWI8RkuOSTTCo
OoKDhmApuDXighcP1tUoquKJ+j6bH3a6nvWIjpQPspXffbZvqgTJMvfr+14aNQih
5/vWoExJQqsHz5IGgoxlFcrJCCExJJV78dii1zJckloRF39O04hOnldQqaxPSFCC
gj9yERLakcg3Npg3axDApMUyPqAUHnVpAAMbDXbft/LEtwRZIpPpSSOdV9Kyw7q9
+4650JkC3cI4I1HkEVJh8n7vjbsoDJY6R3oNthFRISiHo/eM93/VISZdN5gpa65W
qhezjz9LwrhYkPoqNBJhBQ==
`pragma protect end_protected
