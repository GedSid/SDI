// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:36 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mNpZRPknyrFYBMo/9wUtkpIOqRlx1Wn8oLx3coWYUg2VTuULXDj94DzcHWcIb57R
9bG3IAHjclpmpxyGANrgcuQYUpgWjZCdQ3Sl+mwmfIkXMttEq9GwHg32JvkjgBS2
zxHAumeLYenEBGDvmzlxw6aH7IXO5knOXfA7EfHg5/k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12448)
5m0nz3OLWPmFCRd9ZPsr+XQ7pfX94VmzDL3h33Zui/4T1+lswiYp+h9li6gOkTHc
BopYookUhYoCXdgNQMtC7nYQUDAvQg/b3CvVRfgkngsUv9A5KgM5yB01n0CWroJa
3Amkn+cNqbBaCJ+87EAD8BtPddN6fcIaLOsXuYHfzevqkHkKQm5Lx7JFdNafGnsL
cYbHi75EHciIrP4vO/C6lNhv/YnWYId6HU1U7bk7tCaSNz0irPAmPxvtTImCmyhZ
9qkI8ywMjDaKXe9Y9453Je3v30usKqiTO41jabSpr0h+Ft3wCWObwf3AeS91xLpB
8mO2RqAV5gU7vgWU1XBEj1KXaCIpcseVFb9DhJkPYNtLgFFnhi7DZL6BIIeM6egt
+G6rv3L2dODqUSgGinF1eOXuqoMkKwpWYpI3sr7aGfYDlQFMlioOxgJPevwJ75tF
9pDLEnKef+ligiZ8g+mRYFML2XUUjvPWG6VaGyFxIUzH3ZGFLPPONp8Rv5C5hgxn
8DBYZs5R+EiV++rabQjJDyEDi/PjvGOuUIpiQbdKG+OVqyusUgi5NhyUtfU3B0eA
ZvAp7Uyto991AqdJnBsrC5lQdv5l62B8WrqUmmp5a6RP0pIgxq119HjonLQYfEgf
FWAvttH0XXYEraE4fbYmz/Fhkl4va8pacNeZpTuh72/bJloLy7ZQWnzsUL/2aj8e
gGio6SdMnPv0y11B3ROWbVkNq9GQTDhIj8lB4GYkEU5WUt3fNFtWsA49e74Fr7WE
EWBfPh5r3OdAuSnbBPgnOu+YhFh14ViXQiL8YTzb02pJA1rlJ65v2zVPlcPGDIr0
PSfh31vtC7Fp5tA7aw6H/0TABvfNiRkyBI9jkWk0AB7Oell4TjmbkUOO3iYuv7M9
N5xzf6k2Muf0maavHtM4oGUUtuaXM2t+CRI2f639EbOm6rwhtd7Qn2XgXA8r/fEc
wTUI2HagI8XcAcAOmGiIuFe2qL1A3kUZxqgmSgVUYIPE4HIMmzGwtr32DVwZ5pdO
fjVFnFJWM6cy2UtK+JdavUVtDbKqMnq3pZi6VZL+wJxhfjdu9XAjlPp2SszmzSAA
c+SOCaWlHikpbIxLkx9fYnF4HgeiUII5iqImlfyesE4IvrvbGnjuhMR1lT+3T+BR
ZrfLBH952bl8E8p+ADRv/irJVcTDlOac+Gdn/0sra2DiLIXqKgd0U7/Q5JkfZE59
UcLyEPS79TW1PjgD13qG1reQqHmIdbH+1lXKVaBou9S5B1Jw1gWGAZDF5BzWLkCr
apT/H0Zcpuu0LoNZ6CHw8EHn9435w1g8NmEmf6ddvwy/oYXxw9gDTxGhLN5cnS7U
mspM533edRQ28TtUcvRrDaz+l7HpFlnDc+oA5PCPVvtFPBNBl9R+dNM4Hg9PcAql
TeEzN+WCJ4wSihmmFG7/SH6wJhlAkBncRWJUwxmzrYxh/g2gk/wge2eek8QYJcFS
iTf4BrvssMJmC8xurI/HSD3+ddHbRWw0HRdE7CU63zsy0LMcbTpCOyQMHvNryzlL
U0c+kATUWuOmw7PnliCQ2HebQbkU2B/EZAl8kHdYE4UDmPxzaEb+4Ekb8XTckl9N
vPh3eD2ZONRKj4fkSM7+qjIgPYn+HWZTG3ljcInODoUmWieUk7M6j05/iaovRx2K
HS/SVIv2a3hwtnrw8sWsL66ePSqUGwfy8P6Bh3SRZ0Zxi3uZ0fNcLsuPCq+S26lG
lNY6bqFrQD8MwyMHVfQfuodJQJvkR3ustUVNuJzSH14qeSEFhNiQxhuF325bXw4t
INtIMrojEd6jaApbO6H+V7nB76XPgr5twkF+gY/4YHUma05ccEhr09Mn3xm7UUpe
UfL6+zqFfFoASkf1XNUB4HUdKsE2lx/P//S91JWW4nUhnrsk9ZAmv8sZ0lYLLuUk
Mb796w/rfW4tI8/y8v8M657kXSKEbySMXcu4OoYy5nPDIp6cIGZrJwU+8yfpX9qA
5LKByJ37FmwT83f369od5iNRQ7eigl687QJjRUyGHVUOY3ruXqg8QbkZWgSOLkOd
n8mm0L5dmkzijesKbrLzkLA51RWPYRKhUYTSTlqMXbrm4d8Bfgp32XIh7kJZwNFI
OdtWQDBZC3xsiYdXg94bDGZLISA6MoopDKywLf1noFpGKmYCy5oYlBLYJ5rWWOEp
OAW2mrbh3xYaKYC2a5RpL8g2067njJTTk1a81WL6UEk2rj7Gtyur98xsem2RNQx0
HPSsI7hhWeitJXTbUOY6hsmxft4t3ohEnb+J0yEWu6jxJTPnDM8YGQou5ivn4pFT
dgz/iiABxqb7AMwGez/kM8RTDYDHUTil31dqp3Cg66hPscm3dAaDJT0Gi9dP25LV
5LnXQlsQr4AzbKJqbjdTr1JmZzawjnFCP5BTHuoniZwG7mJiGcN72ee7CCKqpJYv
Pc7cRgFZJPF9l4P8Yzhpd4sfR16iC8E2ePEavvHoAeLq4gWyPueRcA570ASOcHsr
e17GYXDflZ6jo3OW6YleOvJM0/qYveBPusSnM31YOD6cVD2i94K+rplE56MtQClM
VuHqmczi1uPTm7kPbbI4uDLNY9x7MyvFTkeMwn+GEfr6bcijlrF4U9F3PQg7nAIF
sn9giEMPty055oNDNbiJ4Ogbtk01ePnFlRBBEeUAoOsTwtqljKsIoBrf4lriI1dI
c51L6EMoXttUCPjEAK2W40hYO05ZkDYgBszk+RAYTKidA/wXAOgPWwf3qotU8ICy
7vy4K3gt8G0un94E79MAjhmVWmKta1mzpp9FYEn/v250GrbTiVU000tEr61tGfrU
Yv+fUwKZDTqIbFoUfatdOWILK+XrqvagmNeFaoA/zotVfElBP6t9hvcbvVeZffxP
d3UMUkG4GoNhCOSVK7nOEx/cnGLCGQrLU8AzeiJY9IGwDV6V1JvN7sIJ6x0Gbo5i
wvug6AcZd9O6nEXQSAXICzPPmLNTxYe7UZm/4zIzGSsy5ACFxX8XEZu1T4KKhq3i
OI8mYWyxMOjdFO+Fo6KP+2xPVs4vOtcZB+wgUR2HE2lDZmrKfsmjrDQpfDMKwEd7
90y04aLHzK7tTA4Pu5g/B8Ksq/FN6HPjNSDhPvUhIt6/ia753AFh93kBEtT4/Ys/
5JEp/oWeKwUh/mSnFkt84KlFszjlZ5JWtnlrnehEqURZ2TXYUQzeFkjRQKPKhAlG
b+U5cHfDE6dbOUmJgz2bTi6zcro7u52sVEEq+sTjkFuDUOsgR0vU8XcQ5mg2WRc6
sJxeGovQQ2iRsx7BDJQPJqPLb3XTKdb/J1KP5Ky7ypPCmdtCX+Wobdlnc06UIBIr
Den2nWBX3xi/0g95roJcNBNcaYh/syIzIreUhulqivn9dmyvFRUiloJJxPSXtIyX
yB8QznyYsC21WE+ADp5GgH1XOsmz7hi7HbTPD2od8L/jyb1nz7y4p8xd96L0BeBr
CTHRsEolMjtTX3o0HRsuOc64t6iSEc27vHaYFyO/kMZzwxueGN38F66AAd1eMi6B
hSAOXsqscG33pAVZninVpXwWksfK4tkxnfBBMo16eL991JX2RXOATppDJ68lmndS
ljow/shXnDaKEM62PSktdYmDKdUh2MIK65CdMFXKlBIZkdsSafxRGcwMOyhXsqCZ
Cb70f7uf0YLL++YWPjLoW5giP4wWeccGElG+ewr32koA3DSTT6KISUn7A/OjxRPl
+WbuuijF/GhkYruV9mNizmuoedL9Hc6qONkPnGJAAz5q7PptiFwEvMZLgMK80ZOY
/2S4VJUzgrTAFpPIANjx/8Vx/VySuRgFv/TigVznh/RKT2VK9z1AdIRPNSrA8o5r
EcodYWnw9qzdLwnedlXAV31At4XvZBHPXNleA59MteThVJqQf4osHB1B88v5pL7O
UMJzSyfWlcjA76yEYbW2az/nCMIhJ1Dy3lYQuXJ97ixBIQjM1jL/dcyokt5r2UFR
sVHjKQ/2bqHU//nRrgOlcomY6+yHHxUzGws5dvcJw/U9fYtxEsdqB4HrNJKyOZ+E
abnzEgMcQogq5fTwRwJktHrr+Lee/BbIlxePU82PH2sbhVh9/UVk0wUIM3l9KRUo
JqsPEJhZ22QGQlmCmtKLSJdLZlx9SQkqVdEIPBTy4KIrMcrxdHhFpOf9fWV01EUK
/9Z6LT+d+TnJEh+RQt2fjrNZ2IAcpdfeHqpXn0VJyJCY7dybM6fonMydmcxgN48l
6vTsZjPpfihZSgWlOW0aBZSn46vjaItDVljtWg9MMtYY38qzEc30O64bbIaav+kk
NkDSbsgoPUEx6sVxf9gtt/lZBbreN+ISNxM7ZU+f/N2R/ZueMjVM+Wd4K3Y4WELr
SpdwNrmVfQI3FG72Xoxy6QB2PKLRd5OTAA9E/t7vbF8Lglv5jU6mkghU5ZnLn9+e
T2v6+SSD7xHaHEL6Qt4ZQHJXvKFMOoOjaP5e7QW7NPIKKfBFFbh2s0lP9aWtuXua
VQerVekVQdLi+KL4ATbUYfGQupsHY0oG/FhWaqGyvjRwfSDh8w/05SApZYiGdbLR
YWXUysUkqcspY6kl2uBQgvpjX5DQtqQXZQ6yitLf5AQ+UXgE0eFa8Jpz37JBPHfl
ewuMBh//dv7D64sIhczWo6QwWCFiC/Oa1orwq6Fyb+M/G5noeFiqVRqjiOIzSve1
lqc2lCe7K1bbMvxocEZy+k9vq/wKApctafKmvjlAWKQbN2l5tUsbyCMBy0Zpp7BI
GPXYm4MARA7l/iFBpUfAuG+MYUen3e1ZlZ8wnR+yX60tbaIIovciOrA+S87BkywU
23d7ccEZVCLC5HP+C5ZA40UBQl5fO6VY58Ua3bFMqEyG+FqckM+Bs3eagySt37Zx
AjmsXpMaLztslXAQJ+tj1QcMKRGTEDG3D49BTKCKxLHEzxiOIdh24OhFl0p1L7jT
o8GjUNcybNIlBGBpKdcMHD8KwjcQdTdpMHp39Nd+AyisopMyapjqLwTXlbIMDTgB
9XIbp/9bC9XJ+sUc9+GV+RFxRSvrlQCqNgU0l9tOoDhIObMZ5mmpIfbzPieC1DVm
o2n+0ejUhDNL4VwsxnM8pbhXWNcMsoOYAXjvWTlgPRBzO5rGNQU/JvZHv06eiwCe
HndPhKLwr3iVCkO7KFei4UuLc5jmW8ojOM3MlcrHTn5Mku7N8YgpRW0hG7QfZCI1
lyj9z694uEoqJtVAEMHrrjD4OOzcPs7MLUpoEFK4iitqSFunBPJcor4lAr9mRHKx
3rJJwFYcRnrXGwRc9TA86o8hfujvc/BuIf4uk7knaE00EFNrkEjC74Ix7AX6zvBE
Tt4zlm8EutTg6GSF2HbJQ5t+go47jip3/FInhFfSnSjC5jpi39EcxtgXlStbwRow
vNnx8R0u3Df0PItOCyA1+fFVWYH7rJniNx4dmgnZCOKaxgQ0tChX3awU+aeEzWHu
ody0BBEYR9IvP96lm+HLdlyB9PRNUsJhjOVAYwXLPe9Zo7QdyMaNBXpWonc+GFv4
uEYCbSGpnEc7k3fWcjPWSDK29ib1Y2sBLX18Z4966Nv8VGYmW3HpywbmnXzYg7l9
2Yvsk+MJDWpyfuFk+yBPYE6URNVFoh++gHxGgpc6n4fb+OTHAw2XtdYfSKhgZ0Jw
NFMIBtAOQnqugDfrhH8GLkc/8fgNTrAn5uLb+gkQDHRJ7/U3ES2gkbGTNofdP868
D0YqcbXtP2xWqSH9R5lQ0SjvJnSazR1ZrUOpEK8Hwr3y9SGq0wjpiff4zd8W3GdK
pRNI8kdfajKLtJXgvrICfkjce528r3Z0gg8yzDUiWtn4YK0NAvGtBNM1BlWWScs2
huNzB2bvzVOjyqjri8MZldaXBqGvpfcC7vA6kJZDXu1ZB/0owRmwa5U+x9bdJ6zi
GWhMHTZzATNBNu9YeVilICw00e+e9PNILRoVYTC7EdkfKevHqjPhJUzPppzz4BEp
gqCwsjbXTlgJelrNaN1zCwJJCDTPUdb3YGW5MQtCa2GXtX0F67GXHE5un6WP0I/K
VbgJXMqzCIdk9yDC2jrOjmL/nTNzQ8rXhoKiGsi6gH0mtNcLyp1GTT6WVCAFQPvJ
+0eo/zr5dCoNhgUJy7j/63fB7wvntxVNN/sNaPxcGckcKzywbu3K6/kicNu46yHO
9FHXMEd/RUfEvJUeU5qQYrvZMLH5aPop6phPZb9TVXhlZD8EYUy8yGQmtbp3vMXJ
ZYtVbrYJTEd47ixA7qG9OrzTIbmu1O5ofh/DAaDndBbe14KD8Gt3vUtI8Z5Zgyc7
ioyOLvLu6qGj+ZKvLHE05aU/Mg8RDzgHU/K6/+xuXHetBDBQVBLbiXy52j4J3clG
XlMwXPnC2ysGoSz+caTRc3AkV6Tcs4LDwxW+phJQTk5fAVuFoFcjkrYpM5eB2Wfm
1JigLbedeWg4jHopRMOa+VFIy+PLzRpqCcfA3Pe1ZWGJ4183GtwkyCaf8PdOQShi
TK/k3L2Ern0E9HrV3qkU5zhUwjjrfzraH0XDMk+JnIxh+YBy17Pszydp/SAlqvhJ
KFKJsG3QJJmMsEivsYCZG55+CGV9XQeeDJhtnQEkmUjcb7kVZIT5oidSJdJx4Fb+
MW3unZY3Grze7DCIpKyVJfpCEePUmzhlO8wLLstAjP4NUq8p0GrtkfDd4WNtKcKd
i/RsGawYciMURD5oy25OzEnTgiPjlKbDh6ydSx3mp6kKDf7GW3x4AwAqgrA0yPmB
nASqpViO+1l+Eghuw3kHnz4IG6gqwnFJT9YpEQc9SOd/n2j5p/6//eM9BWr2f2zv
cCtEXlhzfqgxzT6lx+PEMoWuGVY03OMthXuCN7gPNhV2RXWm9yyNt+BoGUpzIP0m
PDG/DTJlIVzJVVho6BhUdYoncERnxaBDJBNg8pJmnFS83XOvQHF9zyWGCqNXBzEr
ztvekhL61vSZcInxsE1XpDNsexsg2SE5lSdo7Y2IPAMDPp3IDVHJKXv1Rs6W9DHv
Y87ASkhSrsw/FKgIKw+3mBuZ+vo/I/m1fYLxk5neQGm01CS1fro8T30gsY79bi5K
D3Z6oCiY9zaR2gKmWGOSu7Cj4fJdB6HNkgNnJVhQvaQfgqwk5zW34/qHFmCTNQ57
DBSeARiIGJkO20D5nY14VAc/sbYCgoVl9P8SKnxdhA0VL7fxufvwwioS8rtNFk4p
DDo72FK7aKzExGtDOO3ipALPfWLB0xtdeD89VH8bRJNfmgryhmVE6te2N67D3VjC
kciyaddBoTa1kuWD1SNvRttMdo+GMyxQvumeKm/x2ldDj/1aBaiWUc7QOLGN1KV1
XaUhH7gNaxc9FpLtkSYXAzs4oKDquBRfWElhlkJgqkTP3dkpfN9VHzLaGhG11rUx
S4/rQUhS0NuJmAkAEAW5c4twvEt5UK/I5Q64oTyqB+TF79zDS5q7o6a3pYYsuGGx
uJk+RdYYDwsmI6zfRdhWY8t3vsSgsfqNpJJyk/1knneyvWxa/qCkT9pOi9dFRih5
P3JABG2ZlG3iD6dc7HzONReSTwKf9rRDVtkcxTpzr/xPlLVMgRrHYPZpMF0FtuZp
49oW8VJaP0LOBU4JFXRQ1KSCHdhWUXJdt+RtHAeSecDbj9RfRe42D1Csly3qkU77
rbEZofe0nRxv0nx4e3WuAnfHVFnYMdyB+GM8OOLwTaOkLjA2MurtXyAeBLYWb4Dz
ioofSHNVzIm9PihprYzHf3ofOYvL+FjFKep5DHkXM01XiN5vUc3btZamsZfgmJQo
Atu93aZi3sErmfJksw1nR1HCAw4e4HpWKJuZy5xRge18tIo7Q9n5FoyIKll9iN1S
WwxHO0wreQrY5x1V+vXqBUyM0iWn8Yc29/YZcUOflBiMlbBScN8dhHK5h/U04PFy
daqtVr2UPXIVu+TNb2pZbVEPOCnNlAY72C8zOyCHYcvjyVCbB2L8uX+F41lPGjLB
3ytXmzcUCIcForTI/eIx8GnPxWgk8EN9dyXTLINqHrbHBiGoGcxxVWc5yEiO+yXH
5ZBurM+2UH4nw3vCNHnFT4pWlBy3hOX1Q1Dl53HkJ1MnYIB0xYwrqU8257c1iz/2
ZFwDkuyW66ffX7gP9cMwgtz4Yzmor+hZo74SvsB/j2fBGtxsoEboZWzbIryFn0XC
NCvD46lx3bUqIEzTxhRxw0/ZOwy+nzC0X7LSiCo+MjBY4fLy9RnyBDBlNtmRaoBt
G3qIp4dRCsJpr0bCvYp+7Vfvr/zwJaaZ5LL+rKe26ErdCdfWAoOQOo1Mz5yUqMMz
onNOiR+VIDWfZcw2X7k5UmNk/7SX4/l37hItBRMWmu/T/p0woo3MX/eR3be4uvjo
blvRclu6Ia/hOvaz/jXes8+/pCxgWhIx2TLitPnCbJoPATdGAqylg32Y2ichubBK
7V5xAU0IYo4FOzXIkOC/5fx88CUc4NlZypoEKRqW4uRejvPQXrTxRxdFcQtdm1jW
YtuQ3ANDFlUh2Rx7I31hjh/VfX8b/ub8tPCyN1kqVUJY4hA9fzMbSHvmmb8ANnIT
8fDe94MnLEJkDy9OGweFmbROAlTLl0QGpPaaw9PPmVYeOHPHWzMA+V8a63xibYhV
SDl9VYXnUVUW3aq2X3ONkST7+NLJxCOdxn56JerT0xu571qlNkcI3hiDjAXP7ErX
vuB2XiYNVMRkdheKHzJv4377M5Z4NALrzF4aIOp5KX82b80ceOF8LfWcKBv7QcrU
yxszZE8BOs9m4lyc2/trhLOyXiSNTtQ6PxCcaGA76f5p5+/rVfRJI6f6mMx1dvnG
gxkCtqE3OWFpOoMkrJEL0SVuXxmk9UXdD63roQCus2JyKLrRF01eLHC5yvszgXVZ
hUFQ/2xndtvP8qkMUbBOLqiLKKc+S08ovq2B500jU0zG+BWoJY/CStIY3W/Z2v00
4LyXJ3WIdV3JxKLuYaRv2YTjso/W3XAo+wu/y+/Vd8A86BSZg1eFBjo3aHfo0rUo
6ZTy1SqgP0/wtbFLuhmOqULwvqhIQ+oH18oysju5k/PkVRyZXctHMjhzWJ4k7cOq
LCFrLKE727cFNV4jPZNiazVvgNuSxZBeWbbRFJvcyq0VQNUL+cy3Dg/zX/4VCfCf
kuEa2Tj8non/JVeBVb3R2Vsd3WGZtnG14B5Kd0YuvPiGLUHt06fcU+zglKh1jCGj
QGJzVHDsF44Wrtsj3KsNPT51ED2zn9jECkifUr+bwlBOdypiwv4zYwRGYrLs+68d
NmIJa0+jrSRLjwK1rp5eGjMH49AhASvNj7AMjIxj4QGDPuVoy+2F1V7x8JODnc1D
U4VcBmK3u8WhQbF/kqZl9Q6Nq/y6GVfmMFfFwkBicU1OV70EAGIdR38dMmB3npeK
nxbzzhxHYgEX5LaDcXk0t9zkUvlRZoWJdlQOeLKUOKdtsXJOuJh0nOIeyOILNOMm
vzg9ZXSSfwm6hxTXX/CCWcI+WMJZc/0hSbhed4jIjqYYLg9IAcHIw3uZb9mdi1Eu
x5kR3nCrf5Nwivmiu1jy3Fq1BkM2UgWpBz5xYPja49G6rTB5oPJDbBbUokt0cwCe
/Q5j9mpgYWWaKR9lWCi2I47VfV5qII0wQQlglyukILmrXkqttmdDu4Z3+9QadpNu
s1qN9KeYR04ooIMeukvc2j5d9NYWDqga91dYNgGMcB1Mvj/Mc/r/pdefpoW/UwhG
ZM7TSnHkEasFL2DrCvXU0w+X1RzyRYaEbQrCijRui0zR23QrQ2vPBfvbOCBEq5cc
I5eZa3R4FT+gUyGIA+itR1DnpPmjNTtb2cKjsJkF5bNXHpDXvpJTAW0hQx13NreA
uiImNu5VcvTCXJlaqLqqrGPqfZ8pp3fzN0n0X5te/QL43H+EYqPcSLVv4Ue6M7Za
ju+KSZEf9KwB41Yohl9zcWPU78fLeR+qpxc13EBTtaCkGFlL0NqmQzITqAuyXkaN
zOFf+hX76NkYUv1fPeZ+xQtoa8M7Kw5g3JETj4Yv8oilL1tuLNKjTJ7UkprW2reW
T5LhRjC6yjovAqeqMFmbXRHILTpa7Vi53yCuxO3+ieuJgYcmurp3lP8YARJBr08t
NIdJSDpbzLuYwagsqY9w4+PQfZwTKa1g+qXuZ66g0C9p1T8lxffJ0mBNDTC/VoVi
01mGEVGuMD7UYkOeF0xSn2dGuKj9aGRyhHEQAYcGzqn47wa4FJt0Du39i9vcz8Pn
3t3i/oqfdYVHoWjvwt5OH3tnsjSuDDlDelyuItLKQCCpAjhs/66qouXcMxlk9dXN
vmuyIoW03lGj0aAfpcMch/5U2ZIP2qNxVCqEPA5pUhWQUy8gj2Bf29GF3a5+DWVD
HXHf2PQjuJjjkt2p1MXghIBtcsQXBSTAVI4zFsKxMB4iAnaqTriOpJ5+2IBDLGv1
U13g8lDm0wh2QBJfhLY4lsnHImNs8dW8oMPwqHhP+JeZtdfAsr/LyECiV0RnoF4O
0sCCdb+YqzdFLUw4pDK+Jw9SJC+gZ9da0jnVjsCyvKvIeEN7dgDP5iaPpi6gZq33
jlfGLr92YQErTeo/WRJnJz997luG+xph9hSFBsOKUGAo8PbS5EMwgzn9gdNPePyc
fxFI+gmRcwWzjAV/RxIIeSA5JH8AA3/9+9YOYWjfaBhySQnuXFn0XG0CRuPBdT9m
0lPyh+h5YzfYanykrcN/+CdgZewXuQuvUJpP1h6hZ1rRzeNJhxCr71QcoUKVGdXX
yXRw81UqWw2EayFE9+CxOYDFfCcIouoiGCT5cRalRL/NjfeChGDF7TXO6wwef8JX
Kc2ogfTN43wOVdSVXRCu5CB0ew11XgL/OTnGavb+dHgshtLDaccbYSX7qULDhbq/
xJ6uOlvVOTb9oOPiw4MCITuv/cq9ZtR7InVK1k7bUWMCOJaG/bUESnB6NpCk7nST
Hlfri++Ezv32E0YpWpA0s/dW+VFbUgWNEJGBn/GFly9fgXMaT7nMGQrrTUa/sAxJ
nFP6Pq5VmqiwMZeFWQKCwREmIBP2z/Qpa/RKeFJevwtG3+1OrNpJbXAOKBWx2uev
UblMHwgwcQnAtToAQDbBmzZ1P8ItKV7MfmHZuzOcPWdUT+Q3rPaZBiQywj0xycr0
bpB75cfVe4SzHxFLRD++4c4fFwIp6dYIi0/VY2c/pgw5EgOLBx7pnqPaAAUKI5NI
mSvIk81Xdj7NhklfwFPQJOhr0EDSkUpvN4J1of3i2KoI0gB43+48C3r+/WTRUO/b
5ktl41AlWDZRLbXd5snHB1u8kIe6g8eG2/1lpAIs4wqMEX8+R5Fj7YutEP2gG4q6
YbnUUFMh3RBWUFINvh0btOPfA0hr/MGenlvsbv2sdTXAZzxLIXXt/SnQ4Ryo20Fn
Y70/OSiHGuFFqo2tzVXfsUZDMUw40a3soGZ/xCyqmsMcjUb2XBNKIzO2CC/Y8fs5
1dxCfq62Tqp8ERV8H94N3FzxHmiSpz20mPE9KfSK44G2zlV7eOUq0D9sbPvvRgwq
G7V09vwJAYvKQytuj8D9sfUsVV9KmdJd/vaXrHyDT/fnYXwzjj7MHuwkRqaBSqrZ
NpbVIIQ9XZlW1ZLFcPr69Mtaat3Hrc1+n2Qpv8gdodtdsMol9gBSfXrfcc5XQZh1
Bqq8ytHJDxwSrI0Uey+5927+j77GmYhffayVbQAl5aSEogSeVlRO0LuelUQsUspl
SApQvU1tIQFSuGitYwC9/nxDp/V3X67ULYat8GOuyoWL9OWUQy+wnFhLf4s9Mrvt
peQhW/NfKjEKQX46knmIu80dGAhJrbpnRt1aPmNpVcqT78207V76AE5g5E76HrZQ
DrQ3ODUhp35HrAC9dsSyXepKf7O6XX/YIs6BqTseoHTYW2CJtzHfLb6PdYKlAgwf
GfXue+Ea/gzzpEleKX40Xn5ywCh7ZhpybtHp3oBIaOi0VfbCN4HTIQe4DkqZswp7
Jrg2OI+HOHl1EbhJ2q6ZAN5V4iMfFTQ4HXPAD7jrpvxRRroXtC8KxcocTvTPNipC
tYdY0Qnn7UwUA8rauvVHHaiy0/X1mVaxIJTukqiU5NSlE5d5WBfGAj1+P8sAOSc6
wBQY7YQ9DKv0v+jTEWR7bMmB9EHc4WPXxETreCgwKCfTjeti0k6XtEa4FpP54Xk3
qPUYVV9+EncFxJvklwtTWQkMLVk1/WHR8+b6stZ1UhqyTKwjmLkrHnNthpQZPQpY
NmX6Ifke3Lljsvvv/G7vKvhFzriPS2tey+oKwEqjTdyZ5gojv+mr9XxM491gD8Ok
CQ6/yV6L4fpFVQ+hIFYQSNNsaDJh+Pvsgxj0fanU2zvNW9KTJXA0fGGrMOM1e25Q
w082uxSAq75zNBfGxkYN7uet3if7h9F6KJHzrK7YpbgNkCme5xQtv42Dc0MV0Fys
LYaAjVGoAdlj1+GGp0Qz8UeP/l5OBzmhIwMMx38DiJOX58QWr2rJmM3OkbHuxajJ
3INM2s7BUnuPqUSDoKWgx405pySQ55CI5XbZ2jPSNn0YcnF3PWZQ8N1T2lepokN3
6xSktOXfRh4tHFVhta/2p0yenYwA/e0IzSA0LSGXLLQRKTdx6ug+MYHDcZZXPG57
M3WMf1OKoc0/zTsZBhfqfozp5wMwb3pImT2dRxjbFS7LSOvyT7myMWetojXWuC6j
WEFGCiR61FUmdtPGopvi7+w0pr1/Ux/BoEHARiZS2k4tqfIMWeawzIWKZxso5bbE
1v2rtiufgcsG9GXpBdj+We5J4onUV1chrb9qFq9v9XdbvntS3ys1TwsvDn4Ied9K
2awZIco4REGdcUEj2R3Sfq8gN1UwpeitL+1xRWE3nKpC8rmZUMqbeGrIkiDCz6as
qWA4x8GcMaDzVbX0QKOMdwOBEqF0p+cHuMy6GTpKTjgRbMEtHcfQi0nE8QdhKNv9
L1z4VCpmYZQQSyjihS4GjOvHW6OFQCIw537k0FbZT1d1yKY/UslmovSbN4+1qpER
WL0Fb1h4AU9yVcYBQG8IrXfigrfXpNRaUtiknChkgiiQlcMO8Q7VxOQhQ6d/FGGv
pV1J8tRN0OfYXwUeE25/N8F4I2eNWE2aGHUYSlNMN+awEvIys4IKB3bGk6zh5795
qy+HPB7nDeqDuzqnrMzQzWb6Y5PLnHTLGBV+wZyfuyEGXpPXoIj15Q5n+e3Bi2Un
6g6KYH3CKJoj3VS+Rw7etNz0k7DQy4A08yaFCDwiYmHE0Z7/w8oydT2z8eKeF+Fj
CfPSO/8QHlo07pAKf3OOiw+TAtD/XhgSe3aFDncapJvvrAkS0jjgGnMuyewpF8ZV
+PuQYiJL/h1ytlw6s95Qivs/n88rTwnCPy11oHRxBsHRN5Pi+DAsMpOc13/r4cdM
zp6nDqlLS795FrDjelWC3W6NptDWAPoXN5zgS53AOS1bF78IxZMMdHQXEomn927t
Fl4S+npwMTuhku0kKOVNEkt6FfbujhfP2eEPIBhZxLlM0Q65VO6ZrZKUd2rJD0An
0i09oW2ac0PNVMhcoK61vrGNTl2UMVePP4h59WREQXA4Dt6LQL1u4zKruGY6gyBZ
1XV0ZmTCqE0/sEzZYfWysMOxOJhIbaHUhMFeb8P0ep1WAwD62rH31K6ST1tFQKNJ
NMLtpTY+2GMRf+wxPmAre0f1OneJPNq6gTI4px3UYfDnJeIMNj/F8tNnBiW4ecCC
VjvidMwZeok7c1CMuRBYGUiPVwDA5x70uiBFRckdjds5oEWzaR3+4ItNztxJaveI
YpKF+QnGU2qPBp3TdHtzyq7HnjiHOlc+pnJKT3l+q7rV+wTYmbCghp3voopwu7Qx
X+qzice25ABbmckk3+gAvRj3bX5up7N+YTj9BEvuA+6YzepmgI4ksazYgY2e1lv+
YN6huqhLBAaDPYrYuWuY5eMSFvDz2kSWvg2sh1ppQHwQR+EscuPN9s3wEyfJeb44
WPMYxvUQ2JYJR8Z3gH8pNOepGvDDiUzfZc17ig+CkL4rbWIxN5JG12+KbJB1XkMu
lQHqR19P8fvPy0FdQ1XZlA0Mfzn9kvRLjXkRGmHiBreYKFc4lxI8lzyTjSRD5tyu
FYnTvPQFYsWQnV7Ui484hkxJFvklUC0SIK9CW4ndFZRBPLQlZoNK1SakNlW8POuU
1+B/TpWXlceF2qlvFi3HuJXLTSOIyp8ddY3e0UogjnXBHklzKScin8gBNeV7vn2R
T2H2821oG5TN6dUsF+T+LwaZl0lO0DBERHqhiJND3vWTeBKU7QviOrK+2vXMBbdf
fEvLRKz/D/HK35ankAF7IjZWQuVNToSEpDDsTJYYljBtjRtpAwQfJTBiFCkNKtqk
cNSxFlJ3g6NyCC3pF82QGR9VusEeuQpNv4t+YXinrsw2cP+3ox/JqaieCpSXTDhq
MnPuroktodItYhN0dWKro8hLSdv1/niAbkD+jfKXPgzABq5p+rQTda3I7NDI3CDH
JMkB0kCg6FO1KAKBkn6aOqMd91PBFzvuXvvDNLbuBQQiEJJl6aZQdco9Ps+Vr0R+
bBRyl6yyiabkC4Qu2zctMSbaVSaJankKDKL5KMYvVOkPb2CnYIAXDlIiIEzP23zU
+G1sjpE3aFC/Wjng0/hHUI85RX7tUaO3E8MzzwqSfXyyJg8UZJwKwbTVxE34zrSR
cK+aNEKI1tCnKzHI3NDcawbPpvqbW4AlP5UkYWAMJilz5KIGN/ruzFmRUXfgBP+C
/xWRBcsqze8K2piAnh7gtrLdzZDYHm3IS4y+eLCT1vrC3SOXC03pie+4u1aOjB2c
AJe4cQ061qwbQE6zZi7LdmFo/uiOVBTMhhX6Y9gj9qtYCCtJ85SiKwbr0YkAzRFY
440igFqbQpufJvNNwR1JA9bUUC0ctFUxQRn4cKS8G29kmxKJus4pScw4xV8oXOwy
U2yed2ZgYgNrC/E0m53ULhlja/L4zhMcerXAZ7EHPRL7SXp+X1hzXLTlyST2eU8R
LgkI+JBkSHiD5oHhLiumUH9nTiS4d5ZPd0nSxwP1D8m17OjdDvEbRQyF/dLwoNp8
Y+yQZp32snNG3klu/h97ADjAB5G5h1YnM1UQaW07tSrj8IJ8y/eDakKYH6NtAbaV
EBQszIPuSTnm/YrmAVUyobDTjwXCbJ7XsTAq2AtuSG0YeAAvuxpheRj76YPlx3ln
10E5/Zua2aHAGKtKNSghIZMaAtYmDn2/lYTRakhNdxAGDneYOKxI595YUoMRWSPD
sW/W7tmjEEzA0Tp9DiQQOXO7a0RmnQKCOcdretUsAYxNXFs7EldrMEYM34ouNvwL
nVrSgFi+AvVuQfJSsbvB0iMYdq+x3o1KylDfepdf9nn4OaP2QLdQKonbxjL0MkFN
oHXi4P19TKV9MywMAL3auYl4YaU2OLYta4XsZ3xTR1tX0qnXYCo1CMh/64xTlCvf
+5TdAF9iwkpoF8DlrP5skKcXuguMlMvBzXBeZ8UYyoWKuMq8EFe3cFtlRkfbwbRN
lT6wb7njlksBIlWCst0rMs8+zsJUwH3adRrEGW7XeCREwPB33hGhF2rkXmzf6W3g
Umq/GMzW2ZgX+rwQWt/K0lByJP7jTPRgu6PzUn551G/HaETzi98Yvx9LSvEZUuGd
l8Amd/50s5b1reYH6NPIl61R8LaTnREcUfE3gZOBNenCmhrOwOMiUiHcmSFq1fPw
7bJWPlJotCaRreLpIh///yCVhzN7WIWqTlHGT6ALwgGjJq8/8SVU1UWjCaqt2vJN
lUSfIW7EEyC9vqjt96bYGJdzVRu8087/LEYovqJ8qx1ES0OgMRPKBFEa9Gh2UZ4K
nLNVMLYrQ3uCq3q40o5++zMxSmeTBa+SzyDjWs+h2IWAf6QPgdXzonxSHi4agzoD
mQB6FHu5IKS5wGVafTkVLCZeYV4u1orAdqheysXm7Dxl83efcHFUhtKLoh1qsOnF
3O9YaTsnXzUkhNmN55/MS7KAnTAMcs14PAViiOW+9t5X0flprtndOV3HQnhS83t1
jTcLleynvFBmxmMu1lf1M+GDVKCJcyDnBUcnolgAj7a5jqesXJlPsNJrgFTHyf2P
zdE9U15Vf6YSzlUHkqLFmYK+m0B1BFmYdY3Yic/3QcTKzV5szy4+vhOpaBioPI+O
qzMcCvn+Fjd9vqtK2vl68aHz/phI7I1UDvKYlzrMj9Mi2akBQpXuDsD1EzRJlwcF
utgaJjoxhGuNRfTNRAHhfHZdretl4ajvZzcDJ0hXLgrQMhx6lK050CjMvrssFiBO
Qi2txpEBhfe6jzu8Xgc5BMkH2LQeUhx97TB3Xu28f026D/O4oFSG4+qr2Dy/PwJ2
3l3I+653SlxTpL3PZHtZ6g3dAZkvIlVzFocmMXe6XVwcZ8gOOayyvPAcX6YwewF9
krBWtx173fvo4+nTsuSnc+OpTu6eNNuTpkazzPBRaY2P8MS/giKApDOWBlYQTFdD
fT4/PxXAKX7QmCLxPDUxAIUNYSLWVbEv60om8w6i8SBP8K44Z/2dYvja+AzwF068
KU26zXJ2para1cTIyvymRC9V4KKbNEbXn/d6eNvj/x5FbtQAyyzUrVHC0TchmZQx
miPvaOV0zeSUhL/yHe0mff1V3fNRjTBWkLinjNA2OlEyQIWxdMBahhrUoPno7fKT
VDt1piXwxU8h0t3WvyhN7w==
`pragma protect end_protected
