// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:43 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HV5dxLpaN5HTpbwlN1NX0umBQABZoU4p/rRmNfZnNv//TLpkd1UXJ15UKke5UxRV
6Xn0YPbETnRixd1azl+oYcwoslRJbYGZs0hcspW4w8QU430nY8Yhsuoelo97rpYg
PrjogSYF+aU35zPgNoOqM9dWwGzRgXU5aJAVClsKJ0s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
dxBS8JY3n5DgiX/3URpfF4ZMsb8Mm4G3bzFhXIBV/yNaAgl73EVdALA8oNyoLgYa
I/zeLzSzRO+1sQihznB2J/RTOdtrd/ozCMQLzLENkh6/8z23ctc7ClGrSJdKnNwS
vXdcDQNkeQsoDn9i53S5VmEXe604/4Sm/xyE0cnoy3Q4wfutZYePIWu4UJ+qjH0X
6y35IMeynu29UkPMZyftnddv5RQvbbt6pyVJG5Tu9+jRdyW1wq5vUOKSqG0G+RxE
PrjZsS1MicgnajFGNnGNx0dfZjyj5QVnbZ2Ad7Rum8VA15Mof/RU92VWDXznG4uo
ncBQhnm3CXKr+OaH/9/49aHSts44z6bqsalzf1gaNAUJBqoTn+EQITl2yKlWg8ex
2pt1OTm8MXN7hD4f0C/RYaDWSFQskAQzHM0fQcfBwEGDkchhqyeeesypfyuiB76D
gb6Iyq967E2oR6X33b5qWdwU4N3lL3jwn6yBqXQVUoOX8Z0td7qoAYF5M/rXsjVo
v6hSAg/n808VnmOXT6LGjQ3qhtI7q3FSyW429veByBEOqzouL8zrqJJldu/Urp7B
jh1/SPgK63RTiuJ4skl9PAmZIN8AZQfRVYhiCzFCioFs1D7GhBYKaMcyHDYoLEqA
rStmSHGp/Mz83mfyZLjxRx9hzzsqgDK3v7Enqxrw7lTBTJa4UfziSyOY2AsNf4IY
6yvDVxex7fM0Kx8XLPr0+09wihSSULjL260nDt8WEZHypLTI2H/mt/odpozW/hPk
R3zFb34yChWeIUCWujCvREN35+j5E0xWRfshdI16i79sOVFN3n81oDycgml6KB85
c7mjE+JAT8FNvMQZpt4lOLb0hAonIm40GiFT0z5F4Q+F3Kh7Y0d81wut4E4yO+rf
Hm/BmJ6PjphdGlMrA7pUIqdSlUvDj0l9wJBF8ANZNrfZ/lEHDdAcwKPz2HT1Z7jX
/whRWRMgs4E/fHMFTnj5De8QROi1kkXLfDo+PkPIbg5Yg5XsjjRQc6oBl6J9eVvl
fPV8WTZisDdN/h/7Vzn6mhN+CjkDQOyEk5idRGUjaBChCEmk4gvPMg751AL8CCXh
XP+NtGFLA5fjWmG05YnsF7Xn3itpWeO84Q3kVKr5j2dyQw4mvKjLc1s9ewctwR+8
/0mgLN4CCVapN9rzK9/ZwZXXj9po4+C1WGVWBe3uHrGeVHsFPuowSxD1lPYx1uGj
sZdodRUO9v5Hx9v8JhKv/75x5Q5olRpf3sdMxyJtMBAewM+u3W04J8GU6RdiDQgV
BE2WZ7F6wtCThaFT6drlFMWX6rR5T4i9yIKbglsZTuGfiWjUPF9wkt97bwCT9Mwm
8SUGgEHZOWpMTocYJBbTQAgs2sXQcCM0ORfUQtyD+hoEUCCFtW01rgpKMX454bdt
X8QlKx1bJ5rZpXaJjnq4nQtlYYoFmXLVUMcc5WEkAVBwBl3fQfQlr75Y2Zw3U7lO
4PuBdAraMO08fgJAEzierwrUU0A2cfuWiObJhCcPEAnSmclCfeqAPXWKpRK7J+nz
c6nFqoMX4lySSafUx7AWgLD4zAm58lzhKyxtLP75OAtFELT2eigGR9bO9cpKyNr2
t9nWVjOVomf0nCWq1R6WLDvXSLKnugU7E3dZY6Khwzh473yVk3CWVqnXuCtLeliX
QRzi+ZhaD+In+kk5baMMJZH7i0hzPP7spT7ED6bWN55OGSsGJY5qzfnma7b8NQdO
8gzzBH/Vt+BR1NKjHnTIK17qYvtZGAygMUauEHBDLx8e4M2qX3eiLgx3ql6skGgw
PHvmDJgG+rQMp9gfg7FrHXIkb2SabvadHGhguvdV7YZJVCZ4e1cCLbWOI6VF4X6J
UXlxiGNB8iYrKghrqVw5kHUYDnLJlaeLyZRy6ESugG1/FthBGodL7PeCM4VOyMrl
cgB9lTKG7G+xBM0IDrk1BoCW7Whka+3rMXnS2xcCrLkIsXd3KKh03sF6pdx/2Lm2
rjWI6PAZHh3BozrH/wmnTumivcj+HEKltjxm1lhMvnj+DpEkjOfpuE+mIL6LUOHH
mvZ4VDJY6W1AhfMk7BTD63E0RMXSM9+jyY0A2skIIiLImIFa+4O8R5d/G+28gm8A
hQWg2IyGhy1qkOcsv5zIxh6LKHxs4rlaHWOckY3FR85qhbsjSr1+tVH6mCjn0uHp
7v0EbScSvIAIIj5ShnC9o7+LUu1qWiEW96yJkGoborkKWupAnCYLsAK4ZZHD+LxN
OCSuWr9ujhS/JGXlqNQOp8N42Jmhs4NsPK5WTZHDhNl4wGmBLtwbwyWKMr8qDVFM
fkuOSjcCZQexPYnimIJRbtNCNfvcvvFhGuojuPeviwVqdr3eySLN0PxIXi3sxImS
hK5E3JHX6WWCkaeAGi4bdqgAzW4AyGiE6LnmYgILIz4ojwXd0SzZlqq9P/f9OgRo
WmiN7/mQ1q4COWqJmdINYlBlkRA0LTGShTaNEjJrtFZmgmZznBS+aUQ2C1h705hC
cqs4JWAmNVoQ41FPyBww2i1k6khfjLcLQ7p1yxmTwCdgPtBzu9IGwDEPGAQ4020g
C3x9DlQg0vw67Fs4AsMltihZnVOJS07NFg/bHoGoe/FWNo3eajBSQkcGxpzneRWZ
Fabe1UybhBSzXBhDaHGtdRc0028c91nSNnWd1u3o/OHwCadIbLlBBxPOCKorHNEl
Mv7zDaRgUTTVMSmHoVDEWAr31C76qSv+CW2yIgSnNQvuWP30IrKIYbAjXBpXUU+L
TkTWbpXJxkzpWTjClHKGFOnzMHd7vzYopKNnJMs+To8d/fiWFXRkeU3GFiQtXbKB
GzYPUJWgFTsTpigIX/nBur23AtlQzUsyj1hgqmR9a0/NLDPZFRWh4qoj10Q7XBDT
yGdN1WKV5/dXLbwtZaGo2KGmUUAC56KWcJicaZTDav7qKXnC2yn7J5YsMdAWU2Ri
MorgZdc/vX1Qi8kdmg+yxSHuXRFZi/lw2ZUrJcAU4PsIcSZvvIBPS5J6T7UfaZiU
W1HTqz+IzXnRSiEGBGYrhxJcMLSwhvjsD6OeCJLMxdN/CPKBWd4CRfK3xg1CX6W2
etlABjLnXKQTOwIS78WAr/Vas6MMtqSfVJc8u/QehAjp47ZnJjX6IEunrivtOFaF
Q7sEhz/itkff+l+vfGAmol1JXiZwl08GE18uYGN4fXQoULtrttc6lQ1RB2K2Y7cy
BT5xTqCWM1j2uQxErt6Bz/RgzueS6OMjgFhrycjg3QPeUzCsU9jLVMK3NQz6Fnfa
mwsFo/1MBtGcdrN0xQ+B38gLtZ45OaPK6ZKT4MRIaOW3erjWbSe1d0+6w2Lh7IvT
fzPTAxn9B0zUMVsiuxh83he1JbJi2cxcYeu7+jjqNRwuy3jAVIeaaJ4jEqf2pIEJ
H9e9co6hnf9887FoAGM/Nt0/2O+Hj1GiHqkfaPPSKeDdhUj0eBwzCPf6eIrm0ye1
AThAbq7IBwpdD6OC3o6UQ2gi5+OJ7WZNiJxm+EQPMXeP2pcrAowBsMsPfuDNEKvv
PY1GilZ9wMG/j2rYXy9ztIwMSthawTt4/9wKnXdkprTQy5hG/iurd3PKxEr6eYBJ
3TmhGTaUnKWH/HXBsBx6PBqQ6lJoTmOLH89vhl/vDcXOhTkatNftUREP+yDdI5ZW
UZRHIqGnrQlo38FnWa70EeJmwHCHlE8UvuTt+mueoKsXtsQ2E0BYtQ3XUcSr7bdt
R4OM+gfcDBkmsdvC6UPdBjq1RUk6u/uOddwqMpx4lnlzoKCKpNutLAtPb5FCUmAF
aV2X+QMHmNGzZ0Fc66GEqtnO9zUi+qtxcrMh44oWfmxVDha3HyzaMgGFnUPiAbKP
WgARubPoZ+n8ic1RWmSG9EkcRqX4zTUPbnXAcKKJsWs5lOQPm+HVELQZ8CoNcMa4
UnDn8n9cB/zIg4JV7wZJDqR6FD3t3oX8vCyonLUI75ljKmq2vfof4Ll+OQc3LuU9
waB4clyZZg72AIA8y13pOLOJfsq3C5rvY/T5SxMAuBNzssk0qO11/8zFZSybsvdA
37Zi8K0MguNvKnTA8ns3KA==
`pragma protect end_protected
