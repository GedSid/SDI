// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:37 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
su4LgW2Rt6pfxaSi8uj3t3tVf9P2ZjiMIidHM2tpJilv0mjhSLTysbPbSImlPuf4
yZliffMP2bOccRJ4CYF4W+9IOXvQ3RhnUNa7zm548sUasnZefgiHEbfRPdZ6vmky
Qa9PFM3iBCipDgKqbBFsAfbOU6VdJvUtqa/mi3VZ2y0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57760)
oAm4n8BXE1KG3F3gplGnL7i+G8wfoM/ZbtLpMTQDJlF68AEFIb69wCHYEhQJ9/Ty
2BLpnUTKT9l3bYnExmNFR6anGoXPLeQMK6asnILSLeoTy93HK04fIW1gN6fd3oD4
PIgjwHZ7j1+yORkHdxRbMS131yd3W3IKcdiq/zaDMJB70ABoOVtQpyhfBgQhtJsE
usMMtr0vDj4coP17ho/anXlAMqAyTwYvZoIuCLFAsKsWVWvLyOGYJqxtbso8BqCw
y3nNlH430BIhYKZx1BrzYiE+pX40T5eWZuGOSBTCztOCnzY9IPP+/q7KgcEnwrX4
9VaHic0WTNUeHm8xUgOy4d+zJVKuoyfdVwk/oQ74K3n73Sv8GRcag3GFuXNhc/u2
wfS+FD3gUEzjnnczTPR7RcHpyTE8kKMHYKasAR5NpALbwM+5kzKoSkHMyUGRpx4v
gg+/L+zAHmgnr0NZcASh0kfKIxPTT2fHl7yspBUtLbxK0Kxeg8vk9R2grhCXf6b6
pS0a6JNBqtC/jYoOcUKe+NqoazY1Y4gbtRRXeRPn1mSbGBBvNJ0Io3B8shsRlUTI
KKkU4+MvlUfHhfFbPCZCGDCs+k4qPohjwhHp97C/ntDTIfnuYBO5pHOj6QkrG4JF
oJqDLuoitUqoBHmG7P/AQGdcak+/kcJB3uc0vkH8gOetG129bEnCh/v3Z4F2z1TS
+nrw8M5w6T/6wjctB9Ir2kUBQxH4T+2TLSarQrJGMNA58kdoUcU1NWV2s0P5bFsS
U2uBmMQbO0lQIPJ/87pqOA4QXwfb0wq0d074+yoZsSqm+ANogE7I3/lx+QBIyCz8
yZySJaX6cHKMwy1QSqBQOIFytiZWbEyuz5USZDb2h+7n5k2Zjjh1PANNI+5Jqqvw
PUxxQeoHoHm9OUBDF+ZWCawWji681sWldyttLA2Fhi9eAuFTKuHa3tjA+a9RcfSr
MX7asOxPEgIxDmPnuPH8M4a1kMyRnSQINQpe8AmgROv1TUfmfQba9gJRwELGH3t7
/yeTVOw/BRoaO8U7zmxBvROnhZpjH8WAD/F2V8jbdJNxM4WNGCiWRgbmyCm1qlrs
Jg+lIWkar0RoGa6vYr0C5Uzp7PfjU52h3Hnl5uqezh2kBAgfr98k9QQ92eGHBLxm
6Z55B0FiahIuPDEMryXpUoRJlDuFqWpI0F3yCgbgmsHawawPx62T+HixFjk084V5
ScAGB6LZLpl2yRXBHnjB1hpfd9TrfsUXJ4VCTrCG1ifzfzjm2/MH1bZQh7+yjdZ4
n7Ybx+iRggqEgO6rV0tjIEuL8sOWvgN9N22Jh5mBCS4dM/MaO/6UObLWt17MWYkY
1MFdafH6fb6HMbL1Ohufveu1okU21wAdoP3igoIecmNzMpB/zMq0GZsUjVgcET+G
SmLXkTeAKm7K6FKcV5v+wMv57WTV/pv/BTiRROP0fwelvfD3LYHiufHQyOH0jpxf
TuZOh7vc+lAgQ81aAZSwxkUJaPwygo7HlblUNmy5ijPzt4BKi5yE4ZwD29txa0Dd
bSELHZybZe9eUOoX40lLCmTeG1NKHy2by1Yx1CNz4nBqKNB01FQ4apWLm0tbGQaf
8Yt/Fue7m7Ta5wJIiIt0Dm0/OaVmHbF1YOf0Mm0GArbOHxc0KiAFUxOgQ9mjikls
gzimMMAxYiFFn5t+Kr7T/4n/WXnas+RBU/5rhak58Fmc8XIVx+czzxcOxjanLQTI
nbWEuzRUtqK4Uvd+baRxjhg+/G6lV5E7ki11zIRcavU5/fMaPJIjqqzZGCtCWTrA
vj+/pJylkkuP8GuPOYKWDSeTwfcJQQJv2UmkL15sENXul9Yb61raMpVDxcKRHfpe
mJGi7V1M91Sx7lqbBck2yrUpuKclpbPbKp3WT2RchLzcg3ZRZlT/TwsQUUkzZOxr
PRAvuqLJH8WLAzxWXMbiDifVtsARsndRcGzNnTDuZaAQKtpKIMzsKQe73IbTaPBa
j50/e4mG7YF9VT5RGOjz6AH+B6FzdBKqn6sZMCSPCQIZDiAdFe7V1p6TWK4oQblm
kXbZwhfGL/5Ex0rl/Y+VxiDF/abex6+jSKhu1sngiScO1acguv85mqHGCawUbjC/
bhykdLJmnOTkNCz4mZVPqw2nlSKFQ40mXohnNGUSpUPaCYd43UsOSE0EYJZBr7xt
MEdEStS//LW6ZCzxYCfdap55R3CBLVrBWNr23GpE72N3pWZMlFwndE2WElpOjoKr
LceSjtE0AFKug+fpInI5UIvMATuZxFWUObZvbN5J8aSFWkyf2YKJjvjXkY0rLw5s
4P7D3N5f5dTqBJ/wdOG2wKkSggDsAUze6Li1CcVxeGsmNYUdg5fqtC/p3W7J4oHu
hqxhVElgO2CatUZb5HAtBhLl2X86JfwHDwPGJwJ8G4UkvqP9m/3bGHpsB4Ayez9r
zVwQWLWXJBCcf5uSlAGPwKeLgVrRObFsKL2QVF5CJ6m5mHQdpUayjjWZx+NGOknp
v7i6iUiKZvN1izjYxETtg/FwblAwSiJeox0gNrzrZ/Is6GYCqtZRHMcYO2eIxMe8
BclNnXjD81U+nZdsZ9qOuivMjgKMk0sd8bJT5WSAUkSa1NwcKa0LuUF6M48np9WQ
gRgPXvde4n7juMxRju4dIbUQyZbY0iny/QBObnonSugC+iSfShXGB/RF2nnG3jBl
vJVmSbt6ZmWa32clNXufDprCTQ5Tvu0GlyeMILsLJPSujS8DESOrDICmQOwSrYwo
7TCiuT0PghjoBlHYBwlcvle65vk8jV09Y+RxYMEF8eKXowtwqDiWi12UDEzLf/1Z
tUysPE+vSU1jG3RvlSRUaVqQpO9ZJnk1X9BICuw1xJt/2pGV8enSjiOKf3EP4b06
QkhepYZ6Ok1JdXCxBB35pjBJ9WU7nphi50gFrH9FDPNBbneM6KE0iXYK7K0oiDsS
/R/ZGmz5ee5EE00InPoeA2RX0Q+rGW5ChoPOEn2k5Bip/SXyT9K1hjBXItKRE3tZ
ENRJ+CP0M7zTsAOqv7zae2/0ss+6UBELWneMEJPhIwvSfmso+SbD5SK52yXyyS4A
wremHTuVz5oUPSHvIN9m5dPqqvAHs9zXl+LCc6FYhWEsffZv++2koFxsklb4ccfN
7Ow1mZLPOMMELa/oxrFRkF5M9GajPGC5h0DjAUNjXF/2Et3gFNmtkFqHkNlBc9Oh
oVhId5gx3YIqxvHdZKKXbIec2wQ9mi5DxHxt5vPN9/+Qwv+3AxIXFbHiZyycr9qC
cYUU5NAkfTBebKCeolDvnxj9ySCtqjyGkYpaiUeeZtokQVNoyrJ/ylsRdBkSghnM
xFNYF5zgmNEtz+8A3OuBd/JC6pa5Q/3qPSgkNPoCyicSbufmiQjc8RRp3R2zuDDX
I1l2GAHsSHFP8i1eDIRQEt/ELB7jVD5o2US9HZqXhtvasfWjUezM03V1qouhVlHh
OLojdLo37TVtshDcsZwBMCxVlh6RWnDF7r6qas9j0uEeZu92dveh1KYfdLPB/5RQ
TQzx6JXfTFwzx2Cp8uyFGLFyr5e32Hbma33l5YXjSPF6uqzc+YQoimXQb48YA6B/
3wCD18/g/eem9YXNgaUfHbffDcYigevWcLHazdH9e8n6ndjHgoF14LuQzKWcUfi1
ohcFSzyocjIwqkZbV1O9EHrrgexNNKARNmv0WMYtXCZWqRk9ZbdjDt0Jbag9I6y2
fGz5iMOe65fl4zT9Xpq2BRo+oXkDTiVdB8ztE13sUIvDLJWXzolxlboEJEDZDDhj
ppfYFYfuttioUi/FfBRXcdmf2BsmBFI7LZeWPgjwEASu+HXEW5cnMJM6MM4oqO0F
4tip1MZUNF+EtgwTIUECJ8EfBRAsChOKOd3wzVcFq17SCyvPugg0/GgoYlrNjbIA
ZjGCr5OJMvqBDfMo+F0AA2t0SEvFGA6CCfe2MPjJp13DGZhLyo+2TWC+HVBwFuJy
MLxBYpr4m2aa5drLoBwKLX1tdmA/KZ8qfuFI1yCmuPWmaN9hVo9WFCCdMFGWKHl7
NSy1PjKF9hINOIjPadKqfoOCwMwZ+cVlFquN1ElBEFVRxNFjSlNnB47HD63lNt28
MHU6BVTU6xc7cg7Cc4Y2PcfG6/LFWgs46RLKWkLp5IzQhPO3uUzhnWhtHjZAgj5C
8ooLxXPONDvCyrHjzNC5LJnEmF8jKXF5CTj51z4rBiSrBNU88XRiY4PvE2SGYT28
D3BItvmATt3ld9+yOYfQuyxNgoEmf03WHMN1g6ZrRsuKoXkgUq4R8B95XsOZZwv/
IgPkkkZA5JlgrmEAXqWygymujhjDIJGYsmNf4oFoulHpbTt21blyXjar4STwnvNj
pBYbtZdrhovKrC/o2k+DIAjybNeOkq4YY0NBEuG5dIeOHpbBggjoCiKh06Z53FFg
yTQ1oIunaT96K984WLPFBgD1T+l9P0wqSAprjv8dAooDH+xmX9iPevoQTNt6j/RZ
fQqpB8V5ntGsuXApZc861PQBouaeHFagxTD7JUPHx25TjVZrWWM/CXI0LAPsYBKI
etjpgR+f4vH1wZALzEoi6m5hSAvPijd3CJqmZvWYz2x9DGOW7VAufb/l7xWh0qmA
CQDCL475SceHzdHb4ytIkHqzvnEb+fDUSlvrYx7YBS40wTraF0CYen3WRmKkOihR
WGlVT0oKIcsVUDNeBkKXe6XzaBhLN1l0QwdCvFrLOmgGoK00MrD0vcGDcVhSUaBe
ccthuolFYQDc346ruU+e/2atK6OEORo9BYX9sTU5c825V+9fyrNkrvtrt0snodnL
A+vhn3J0XEFR9EFnG8fBFFCnABkcVg9Iw1R00Q2zvsMzHG26alMWsnJIjrx8EtjR
J2EzsxD4LLdeP4GzOSPkCp9TNn9W0rKa7AymmF8z85bWOCYrp4pZPuwVzi97O56l
Xd7gZylqmLDWI1DXqFNdEocURwT4bKmfS3lpYlobQyPtJ5JLaWxOnbWc+lXvVQEK
HF4CaobQm70A5aYuQyUgEbJVBoV+GTznpztkWtfcHL3dHXxsPjKxmnKa12Fn3ldz
CqL8oOIJ5AYIbpdXZ6553E1J9H9hIxsrPjt+h1WIfCjQmm4U0vxw6CW3FNiJuVlt
Sp+qT8tQjEX8gpuYBNV6X4X7gNi4tcan+6vwex6QJuEI+OotWTC9OUXhifLgZiP+
C23U2xF+t1eFX5jcOkeo01AtUn6kxlBuB0zG6rFV5LUy9Ezwp8rdkBQiLJcLcjQd
U9YyKo59SDTCHNFNwVTXc/Algk3f1yRc4qKBDsO1hJaa/EOSaz6qSbfpUgrCl0Oh
Ye2rULRVzvOIify4H1i+7+XSPo+gNilN9tu8KjAMJR/7GOTlDzul2cOFy93JF8yr
VtMGmw3+uXz4gkSCd4kfWEvF53fv+iOXxUBbdRBvdKyTVY94y+HNAe9vBuIr+X4n
Jy9Sq3F5M8/QRlppd2BtO4ZhgFAEqbqayoL5lS7XwZ9UnarGXqe4MEttVbNPm9K6
FK+5F4mjYQcCOpks6x+07ZJQEmI4EZXANrMBr0MtA172dLUXGZU+5ydKizCvrKgZ
5SW2pPAJrKemdn+qIxc6alxVuNgpqjZcCs1r8qCyBaq3EsMcIFdVQJ624DRhJ3Jk
3WQJHRscAgtWEVaPK9uLYItwxEEtsdhK2R+EJbPXU/WloURzD9rNPVoqm28iANcR
QNRnp6Vn7M77gmBdVtUwTy+PFnv6CTe5yp5LiXX52i3B5FLx9HOq2Tz9ldCKtP0y
M+cF2GPToO3TgsOnfMzQdVF7+t2kVRR+tF1t9rByjrzABc8vg7a9be8TdSDi0f27
VCW8tRG5rG0EXeZ9izglG/wmNj4R6vKJ5lSJKAWVjP/7SB+y01Yf2yoSh/PUTMfa
7O0x9ZdwbG5ATi31a8Mc3dQpMTuaKbkETLCDZMcL2BXePscQHFoGf6DmAPTelPcW
dCWYeRX1jE4DVbS7w9xOS4lDKri7ElMD4MQqeUxCeFG9cB33R/P5JsVaZdYONBC9
DO4eHvQp6ffxs5pzgWQff3KKd+NWmF95Mo+uKtkprZvl+rLyLTqs/Hs11aA4N/xI
xvkOgKtApDCafGRsL6jdSU6jbHxMiUHFn3ob/FBIt1TJVWzS2ntqVsaXFnosXDCF
w7Zq+fAigjvDP2clgt9NSTs5JSvjeWaUKXPsQgW7Mve8gobYPsEGQyxglu9wC6JH
gnLEgShtpYm+cxdE6x2xeJwD/Jq7YMUL9YSNjMxuHlyqHvt/fxGArEWsU8Alq9Md
N4c2eEmzie8Rei+tm3LbMZENYJuVVeYRhL4By5RGl1PoQhfqc7RQOchZ3OseAfFQ
cFhqaEakxP8Blaj6EPXIDMXOCE35dhrhCkDdzutkv8d5apBBMZUNxLV+T+FHga+D
DRkcdU399N3uCG9AEBST6ulXsCsVcRcav4c+D0Lgi5oIWvMvbJV4o+NIYgjH1gPi
1xRpVjnNAs08t/KkIivajRO6GaJt9X2XAFZS3cfRlibAiuihXTFbBhM10gKsVADa
4gygctRBVh7fwduqZXRL/KmXBqEMilzIsg2NtJ3kEs1FFxUY22bwBJ82IEBW2Qb0
PUb4gl8sJZrbZ3UmKKai46dyPesQV9JGIVJU36VG+s5Th7ANWtEFswR790velX7E
MZbjRmC1IcDIDWfYb2ZjdOYQvzWqbaC+YF7HP2Fyh49Js1IEUUjjx7tlNIRl0c8q
INQkEuBSBST/A+SLt0hApaPceFPvYgHElXHiipuPIQOcF68mlpu+ycgBObLHxKmW
r14RSEGQD3mW/ruCmf483BYb4C/LndMadVv75N7zuvg+doddVI/+YqL15u06D9mA
MiTyliAw+3+AJzQAIQvcD7OgU0178IzUYOCk2B6r4/uAJHZP9sBVzrDh6WX6E0e2
JEB1eaCMFJoWZbD52nNHk09Pa0YqVuuxWZCCd9dukUTmNx4NrPI9/Q6D9bUgKB/C
kO0cXOq768L3Y5izVq/M+keXAqVm6VjBhcemwWF/vdvZ+zXrxEFY2hE2QeeRl0xL
MEFVvYcILUnWO8WBYtLP3mdFJ1RSDp+b/C8WcvzxIVguA6ZmVkFZkp47/X2SSFjT
JsBAX3+xyz9VxJfEOVOF6l7aYKX1SGSqpCvov5YBL8i8BLOVlzDSbYsSA2ckojEM
dBoIXB8tOj81+ucF5pyUjLAKkx421fC5MO5ac8sIyEd7firmuLRwMy4Js9NzFxPX
tBrsrWkfdik2EHxfzSSpv/2DxulLgoBdecydPhkT6sTTSSOVUBTzLf4E3TmOTKyF
ZthZ+Q3wOqkWtH7oOENGUpWw+iseRvJvrZHwNMi+aj3ZfqxwaLRPawaSK3u/KzPj
NPxJaqJ7Nt4woxVTJ4V8hFRbBBV8MpKtSWDSKdkTzo/i58Yt26PVChPykZSONNLO
40Ay8cvaxJYKPbj9KKhYlNnPuvtFEOekOjd0CYo/aKjzdAoxPJ2YVyh3cIok1A2n
g3EdRXC5262Z25HmOCa46CpgSl/LieAGLBYf54vNQqbwZM5zt3z9nOxXqc0HXqlW
wbWNqT26tgsmiBgfj4Tgbrgc64Fcm9TIt7nVcYXOg83AE+PrNJ7Cn2y3u9ZdDAhn
et5uAunTGIPgREsIXaU5cBPiPadn1kput8gI5Bp0580PEolBsq8PVACMRlNvcsB0
bNhmUMnKAJ6VJJiRqK2IsK9F5rDBnyPTQ9lGvSNjBXyvcba8paACQ0fEo1NAikzP
r+N1elH2y5bnPGyAXKgDKQq5dbaH+F3XWmMWAauY/DePpwMrtWR39cvuPXO4LF9J
mEDYCGYTH9igqxgNS1s6u3SChjg3fe81rVAng3CFhsqNUeTQMpzdOJb7m/e7fQzX
a7CDdUi0l/PB700QEblnImL8BufRhNgulqGzTesZVpfYWfcUEp0exnw2EGLlGRi2
ImUWuIv6FECIq/XXwrIuRWYq7hoL7eQCyOc9RZSYD69GVZazJeUMk0ymeIXZa/eT
jbtIRcTUQWqI1AlGqJ9f3I07KtPCZCn8TFOu4Pu6DNFeFx3LWqhFJq7k815TuK49
dEj/mHsc4JK+VvjaJmufEJETZ2AfFWPlBL/AH7CKRgfmlT5+28nWhSrey3hTuP3B
bU9gfc3AtGOcKl4AM5PRZPbwlBWTpqJ5yD3mVvz7o9WNby/NYs0Es6gDbYDM4FBl
IZSGaW9+KciLxM+bzhvX/oCpSXoxq8+Sq0pLmI9xjUN9NACWKGnEbB3nYiltyb4J
rwOrQTeY3JNDH4DK+pbRBJ2CRTFITcI4Kty50sLKL1Z3xZxOT7hGcy6TfNrgngHS
EkRcQ69q32j/k7SM0Z68ycrm3t+t+NXZ+DeaGH43kBw6L8ueN+p2mDUeYAQ8fT67
ZyL27TWzS5M3JHKEHTRLtjpwIAaXEcbudrNmu7/grxSjo6UlEAEc07zjWKJdqK9u
gBSn5yhpXstx2GMX3OcGSe8kvCWgYDZrVtmBIIiEXe6HimDYhn/Ox4mf4eV5k3yj
aDgK5XUNlxG2yJvh9AgaTMQKA9ho0/uW50TYyNpiXgPLuxicxn0P/3krmkrNxj6n
VA/BiYU7Msl5M0BL+Xg2R8wfvzMnYTao+ofPW3WN43i6CG8adI5kxbgE6cI0IktX
ehTygMLwlmsZ4skfS8WlrtC2XExQPKFn0E4c1pmxhiqTu/JHquM8U+s8z6ooOD0o
IuhygpH4UvqEjku5JSMNY4yH3ryXGarh1znWVINJ+Wey2FLURCi5z2TgUmcpZFRJ
WQAeS78Le9foWIkOb3dbaFZoh5SOqfhdpwNmMwj8hdxeAbb1NSLANBVWEBcfOJqo
NrkZS5hQ5jhVzkhdqc2t+Y8+nHmVZV9GcQGqD/rGEBuxuf+RlayDDAPDpJkwnWyq
aMlVE/GHgQYBfk4kOCYvcdXjgo8K5zljAlwplQ6zjk42mRugFRX+6Uv1c4gP4YPj
QJ1nnmq58HAk6+iEb8PvwtpAOJary1MJpoqNNB9d5K3KOl1j4IxDnhsN1bXb+OrX
PxIfdY1irMNI9Jb5UGDJ4/thYlCLHKlwBCuBYBVGE+MkOzUSxcVjWNG2y7kLGpr6
nPH60TDUOvu1DXsOkLPFbZ556hb0KQep8+2DrVbXouz2xCx8kbx915+8lwgVSo0o
GW/WEldqrRBUfZf5E/RfaE98sjS7sE57REu5UmTW7XJaajUeFYBEOfIVxUyMsGMU
8I7J1ihYO7Plj7yqyBzkwcxnoOWEEA7IL25QZ7FcUXiVi4zZwZ+TMqjPwtq0g9gw
fniixHS82fnnRM/1HlZ5ywKHL+OhX6Udx6FVdjSbLO6QnkSrNw5sXzAfKsrU+Crm
npgFPzgAXyK/KL/d7AMP0ElxrlI88hVDehwSWhS1G8EoiL4tsd7TuvatsIUyJ8nC
TyreGdtjbxZBii5+9tqjcD46mDxDBfagdCfvwBSuIZdYliTb3p9FOdajZW0s3TZQ
In6MihgCWU5t0qpH/XEjrXvhfJ/B8B92pKQ8RGJoNqS42M6WxXLr7BHUqlInTHtE
olF4K3T/OLUi7czQ9v3h6U8GeqXrLvf31kpFIeSBAmsQDPmLbN3sqd3q6FhvnPMh
epct3hPkKgsFoELV3eURJFeOJDZsqBHa2sVa+BcDjhHHAidwm1tqAe50PF54VXe2
eABO0WD/2u3KAlaQjsTL2jLtdwqzuwdNPlooJ0YnQp8znvRyZt8thCg4S8sJ4laa
WMPwXjRH04eDxbiuON4sPdQUed4rXr7teIXoXzV5kw8/VbflzipsWm3JZkLqMEmh
tV7ECxM9Yxf1fTBcE6UI+quIdghub9Dw6jLPJFsptlhWREwG3WSf1I+duS7dIDoi
o5MKJ+tg1fpR57s+uhXXYv6U6Am3NtEvattJCY8/IT+mJgz9CJKzm4sAmjknW/T0
kxu9e+cX+GYe6bGjSzZc7RmnuJwOIUThKzo+YufmE7vgCPnJzeY93RH6VVWHVyKE
W4YWxnKdkxx+MIqWGSfGDFYDZZ2TNFlVvtf3ZN6w4VzOTZqUrBYBuNa38im9pqFY
RyyeeU6zOU0CAdmnShPgRhJVNTmyHdOmVi9/uFwkOP9PG+AIpBhwWH0FKA/zP1oo
QKuTAYnoUypNjQPTTWEeafiXhstvsyqRCA+2uhzBuf0N/TYryAx2GVB80UFu/r6q
JCcP9TDPv/VtKAMrmo4c8AcWRmaB9IKdfWcUZwelmpe8krfI7Qni4fIoGLrKHQn8
sdLfLLA9GXzFTcIOMRPqgob7xEjvbaNoMwVu4u6jeiLA/6bMwL/VgZ5g7Go+TySC
jyTtdQ1D8En+K9oBUgIjjjFpyTtTxKhZ/ivWiaBC+MW9QM6obcRhUoMG5YKVxN3g
EAqIhZA0julUio77uow7sv7HU5w3QiBnbO+R6mLQr2ELKhJgssoj+gHnAIHhSROE
ETFT/8nkB1KOS/YzZrZcGa4FBUgGRJMmwZzFGRkbtR4+dNQ9vOST4MofWQE5Zmjp
IFjFVFsgBqecbFk6z9mhsKSTGYKeuQ6MpKwM5qhrU3oF/QduI+NnlRHXPyvm5V6/
kwZgdnpWBmwMOe+9BcE1LmGXMTlsyk2nhj7KTabT+EcDm5V3CiSKVQwGI4MPkjmO
+IkgRBmXJAHpIIrns60jfz7ejAB4oMOeLzMgOgP4Z5KBtKOUWQ9t3PRueEc5Tap+
xCYEvwvJfpBjT9iUTpCckF0e1ngANqF+qNi612JyjjrPUQS3US2h+M3Baw+J5bGv
MP4HlKr0aVLbDE0zrgruASz+WeTMRj/t/NCk0oKZlL3GBnQeSm4HWiFSGuGtJrqF
oVXRtYFHGJlus134m+ngHISlyxZPASL24KzN8dIkX2RulhgA59kK6rC6krGch34P
NR687I7Ek54CetdtVmNqryz+V8PwCpHBdAWDqo2loKTVTmY5bXYOMwgKrQBgEF/z
KAcalnyrNIWwqradu5I5XD6eIq442R1SNNVH/K00Wnvjo3QNOMM/grMO+x1eWc73
Yay4VjrGpth9pbrn5WnfPKt2JdJBwrw209wsCUQyZfOFv/OTRW98fyMsuvHW2acE
FtiYN9QP7Obktc7Uqfcxbo+XcHN15unCuZKEPrGxU16wTy5COF3V3FUSiNPttuEM
GLirMUd9ARnvospS4Mrn0U6GI1Qpu+8kSFv6mhSR7PgcoTOJQsfahac4q4hQurYk
kyfSLzvMxBGhXor3mfGXaHSRsWxE+Ti5D/yL0JbWobseSTxearYRGpx877TbgSU+
g3bHVOdC5HVI+oc540wxBWDbHCNg3o1fp/rXpu1XLFW0hj5VfvGgh0Cow9QFk7YG
d40sK/yRmztKHh2/yNaiGD9X0WxucSPHYFbkvqCahPli9jJAfHTRNvFjsk4igbQM
dVkueVUTkRmQBzRUBa6zm8LxBWbCsqKLuIrpupcNq4s1Dwu8QTRIQYfWcD488cd9
BmA9YKY9H6tyuLs87hcxVYjVqhzIsOQlclfDLMQUp83TAS/XJRZpezxYTwP7EG+T
FguEwSIRoDMNGbHAkBo6zS51ci3JYyBShoIbEj3K4N+MjI/FARUtIWI+udGdH0al
e0Frx0S7irWr6ozoWlAEnYnPx2VTwFtGGxY2oK7vCv30p7T93iVmiikDFebu3xLg
rfhWSCM8SZf8pluj7PNbj+stS/PG7WiOSLE6LYd+hhRvGWSrd27ibaOup/FL++Ea
sApk5yR+eVeegITroi9bbXhmKlGzAvsgpE+xMMLjl4+cafRU6xLeek9tW9UJkPjp
HW440AS3G/9z0xhK7S4a+eZcetIUg442UPberOg2luvEdVh2Hjj5yePTNI+3K7O1
C7NsDcci0kLqCzchbEJev6GmAvnuZj1Ux/SZVdhhX3LmspSRkgjG0v5QiWa0t4Nr
NLa9/cU0yGwjEe0WDQLt4HJQYVrAkg2CYwnR3XL/pyz97bbLuMXQaBnVwxQWV72j
5+xZanVOADL3sJ7+SLJ5mpSh1zi+82Y3/H+NKfaPIPsHguuveZLGLRZH0HhflG14
M4LBH5AwT8BJi/t1PZ3YXGjfJttGtgtfj/gXKgc1V3muL6ZAqXW4xXgGlDKNWo9s
7l6NAG27RLu4J6AuSDO/DY1HnlfQpPD0CQtfSTXN0VwkjcQlA90ajIuth7Rjj/7o
VWXk/B1tQd1j3C457rZi9ti9Z3A3nsXT+QYy26tJYJi2N8CVzEckyFWSKPJ1vieG
gcg98+9ToO0NgabJZ4w6j5/5r/5zYGfdniovRLfqw356NXW2lEWbI30QluskwVzx
Q7ohbo1jX6yG/vC7O+TgYmah2Mw5dZqP3cTGImqKyztSPdCcFYNTj/kqMJJ8tUY5
13/eLvATxKmjBqFbNKhHEtEbNdd7jm7OmcoSvm4h/2sVaZ8aZuQdyoZvnvwWGCrv
zU0FeGxQkBZtgIIgTYzeN3XTT5SgVLHnI2fujt43+2akeTDrXDbDDWix2sq0+RaI
wG2JgwuBi9WdyUE5OWjnmrQjvx/6Ec2VbVgaT9xxabSrZByLk8f/4wTFzfJQTn6T
6zvH+ErNuBs8AdtyeGk46lYXt4GYk4Ne/jDUxYFBWwqqCtMjSoLsVQUjupB8E0g9
TL5o/OSjRUU6CHOzk69pMcRK6jpblbklCTDxyx22onY4sAfNiiby1sLLehTtIaZs
0gyFhZLfjP/r0q13rnR5KXIu13G3hCXSXVlluLY4opYRIGEwmBnwTYpJMnh3uh80
c7On7IiCUxxOJyGsq4QwfSlXj1Y8CeNidbYCtj6NYbTqMn1R7It/KQhgrVVPw2UX
YBV5KB/vGlLxeBne0jv8br3f71RcHYf9H+flNyUw3J8a2tGKUwzu5/9ek3bWf/Rk
6RmcgyTtBEWJwy9RzgtQNgv8MGLx519sfOPjQM3KKKaV70BnTcd7466hFYoTjzHz
X8I5/N1E6JWTpbTYwqLwddGaTYUQRTWOoHzDXA7HorEjtYIK1+QeFfRn2/knvGnS
Fcx4oWvORe5b9sUXZbIiVcFmw2SjpOOlCZjYlJo+eEc99ZIJA89wfUEQeh8IwPaK
bfLqOQNn08jOEbsdeG7VnAdBNAGZNVpqhnQdMAaqupYI5WQoOpNt85vJ7bds1DPa
+G5Kn8+hp1SpHbo+BsVPDJeQMBngYuKf8f1WBjHdLguaB3c+pP1v9FRbbky22L3I
iMlWw5f/+CaEcnGoqO8Fr2HtRNH67QLFx/ZOIf8I2f654qsGvKVLI+tX7bbyloR9
eHIYvoN2FDeJJdfUtuTxTmA78Hm3VVTGQtPRFTEeUugKAYK+Pm3xIfCkaTNDP4FU
VRxb2KXpqMbTLjdbI5IqqdhdtETHhyZfrnYStjj9iNxxhm9ibAInEOixhx3h8ijK
n7kBudlZv2sF/PoAiJsJmG7O7mM/9+w7poR8YuyDSJXUC+rng3o+qmksLeIGQJX/
ReAaq2hk2W5B1bECGbJ4UCDa6zWxJcTTFnepZ2D7w1on7u/5GjtnIvkWs0PpWTxM
oo+W1JPFLLo6mgHAkzL6apMmBJ+dF2CrMqvnVy/E5OCTSIOhLQuukckWg/EE3iHH
glDhKiHPAjonGV2Hm33pEt+6OmfWJefzoRaRHLM1lHfnwz0RPzCIRDO+RW1A9s3x
5CUZ3hjwLemoqIolaD8cgl1ZaO9TDSxI5xWD9Ily4VR6wdp1lW0Y/yUd/lnLl/s/
/X0Mn57kXC2VhFa4Aitt8W/6oREVDmInBaloQpNlx5fF7pDCejasdBKS40WmwypV
Ma6pyTwy27HZTbuDvi8kcyxmfvCeTF/HWdRjo56J9L7RXiFvbSpzFFIPEdUgjc1h
4vB/S5yZ9ih5Afjp1IHQvr3y5XQNDwdr1XYRz3pGQH+HurUGghwKC15vwrCnLGkd
0bjHaRoJDxo87Lai3SgklcgBdmt8oAcPiBwdeFC60KTtKJExDUSnABh2A6ZES0y1
qIKDBeBUUTZoP7hDnMfm/5oQYvELX7vmo8k/NfhgVsTqcCXe+sOYiNs9RrAGSB3N
hxs+fj0ITKukZ3OrUnSqEbNTaYfDo2LdPqxabtKRN1w8uRT6WZZ5rF4p2rBRTadG
d+VegzwRjSkTzvfA/yAniWQkt77mbTnc+ZWRibRl3ZJIWdRVAqLEmtuxYkylNV35
aWYHARgtXMYL9FK4Q3+B+/wKHx7I6Tr56PjOiYCQciaTeCRVoZuoiMpFWencXRPQ
h3HZ/qZFhxgSvJzDTB4NxCwZPjstjYtWYRE6t98hBWJhE2muMAQFe8TSowNGxvu3
qCSo6AfzZ/PlIGEMwhq+Ce7VidfLFJKgYtpTFRbPyiyp0Y6XYkPO0Zts+NDh3Xjq
rB7syAlIaahhOYngZDI5kDBrDwprGDx6m3peYI2g6j4JUSthwoUa+f6JSeVjawvF
oSQsZ90ZOkiSSVfcOxYWCR1cUJExCJQypqR9v2GZTJ455gZPSKPRS3yGcC1iqdws
WHLl/cDsKppYGcFxUr7RPWXfIv38O9y5V7neJH+54fIYlCjrxjKCpk1jbL5/ABq1
yTf/Iu+PUYKE71KkXZH2pY7K330Wy94w7SdHK7nfkDV2ffjcgRT4G+6Do/njCYj2
RnPa4c8LXqtZaE6Vbk+YXnUkQ8LhtpeF19+UYpLHbbfoaYgikXvVuoOOsEVfmr09
/w6Pq/oBcsLQpIjySE7ghTxT2qmnVn6B151zcJz2qE4eSUiyKyTTWfrrW0ZjNGFy
VI88skt6zh7cRgIaK/dk8bepdOuwuVCzXnagLzU8/auOOVwtQgpKv0rsBlIetmo3
VOKjS6wf8+j0cvcICG9t4UY7bMuSYQNnOnntsMZvtqWi871Mas9stmv8Pk+WmjiE
v5KhzcJjoW98u7jymetuPlWeg3WlSclN8y47v/3jSeQX8t0VdhF9pSgbA3jmK6TD
VWg0W7p08m929OUzvSGbO3hy2XD0DVU0FdZ0NcNEKh2z++hYng0pjipbAh2nQQzS
UgM4K9ykFOpSXAiG+EfrB97zDHaX6EH+AUwd0B+L1LbwhIE2rDydb/8is+AEoz7I
kVCRgnTdESoKfXskkllFgvQJJ25hLp1u6LH+y5zgETr+bDJt+RJ4b/VAfKI/s2i7
ZoUuMx1wc6FU1NnWraUEDSYL+lpuHnyW7PnZ5wfB4F6Bz2aGXrT3dedYbgYSQAtQ
o4RWagFtZGdpHcXqE8RcoVS31amwkj8Cy+hNtYZVwao/jHCJ958/IR3cRT9ov3fB
kA0Rp0dnMptRLlPH7X4Ni4TouKndEmDvgtbeCkgVO6Ou+GUHlHW1ThqyZVvvYT6b
4K9W9zDuWhYQxuQ9HMOgoPehDwQE8UC354Ja0PQ7iwtn1Hqrdfrs+uKhYUsCrkw0
f+QkiSC5dgo+/F1hFuhokUT3Zq7doteQ0llXWIC5Co/BWoMd73Jq/duVAkAzoXlA
Bj8dGYeLbSKwrRG4sc/tMBHw8n6/vASYxj7VbImpydPHtoZj5WDgiDhNoyRLa1yh
9yt8OZPhaf9WWSmmRti0wV/Eu+5bWAxQEIvAVaablCYr+MbgRul2ahRi1WNQ+Mll
WcTBQYUXdhPoR8Dtj6/jGSN+x6XXqp28ER30tADWewEJauuCAlpHtQkiIYbIUYtm
7XboFgELW/0L9U8ya6///myB2P062/SdMwa3w4ouVw+6r/70sSIp/GdNL4Mt0FF4
mOClaJcqnJaLbPKT9qMUyq8aMDNuJ5ji2HYrHQJb/wUeOZnjTgJ202Y85ulcT98c
WOXxXf26GBuYnqJ5uPsurOnckKG9s5DrzzNa9ghg2XK0N4BbIdeZ3wmJ4d7BN5dO
CQxZmqRBDJh8G/K/iyOV1tn/2DGueCzD/w1AmNtOTOnD/ru1d3gd/hs3blyXGP8u
2ujxd9RPGh/CnXqGjf70ANUoe4VOCk8sdUbWh3pUhsT0JZq5ddHdhKm4Vn0+v7Co
ejABv10+eNz/EC2kf2qQhM1K2TXZlfB7oE0kHyHYZU4aF/wDonSNpF271m8VFl3E
g/RUyqdZ2EiSdfrJzoYKWJmbTAWbTD2lp4wE218OhuAijo4z4FywaQT4fxpsaf95
NOpJtM9jGGhGeSQTgxE2XJRNETOAbFFaKlxU/zFAwVGb1FbQMZbZt6E04S877GQs
L3kT5Rg7grUY3ydEGWpyuyWc6GcgczC+lcsQtCXdEAo1ZiW7VOnyjKBiVygxB+yW
/gmb824WP4tYOZB/RC2dKe0fOhXj+onxhteiMHE+fQo9vz/r3xr+3063q+tJIJAR
3lOt5qOlB7kJVFP088E/tQzNBTbsrDajzLAnNGJ2f5XdjP6L7zvTzSILzcidPgPv
Bk8GTSHQm+pwh6T0gSSehoZh8Kfnh4cdnT+KqWsD0h+CL5asm+yyVxT2FdU8HJZA
0U4GRrnYfmgOU1cMxaX4/5yq9g3ssI7aoKyOnfe8K+rOzaV+UwBBR+fe7hVpBHLL
02w/ZhIhGCthMzdURsUTfxpa6yXsdYwee5kRaLI9F4L5njiQw68ejJOd+K1ZLx7V
YH0CdtPNjS5syxDLzpGlg+rVfxJK5abpbT46k/f7qVP1uTWN7I8os7IZ5xDAKU44
m3aZUeDVgomLArXaDqoiZ2iImba+YIAVm+5Qz59mXoLb/K0Kcr3YtqdVjaBBb0Mr
ViNdiEeugwGdGYUoeHFM+Mpx2Xup3FrqrcPC0X8/Rn/RHE52HCJTW9UfCJv8S1of
BbD6ru3O0z+lHa1HYx4wwP2s2pT0+YZnPNwNlxiVUbEbTI84b06BUO1+dey9/Fxe
qbGbw8YWyzOg1eRkzWeyvOazeXnfnNe7U/6u1U8QuYFeku3VEDJidqPb8DcRzvHr
st7QUYa2Ow1c3L974l0Tm+zVQ3qJI+j1LCr4A3KK6+jTsD13pVvzvg0/FcY2DN3j
+wzb2pUctWoc/ImHVL20oD38HTuKmzxqQzVeH7eJOGg5gr2Kw1vO2r+wb3Pswe7S
iikFXs4DFZBOTiZnLepPZJ2C84ouPlhtg2yC10/mN/iw9tAS92GHdo98Y+q5iyLE
x9Og7Ke2hd0E4U91b4NWdhLhiA9Hz14JsjYbkgGmL40T/dGSf80VkL3AlrUWEyrm
R1M4IXmzE+YA5hM7ld5j8yWtq+0yWhVEUQ8vVpNp8RXQY4BIysM2LQ65IG77WXiP
jdQPT0NoFTJbWuSnXozSBtIhdYsZ4No6xiNpg38JHuBD1fnKABmZDsO26VSGxTlT
EZCbM4reMN06n6Nm5mnJvfpQXgtd7CcgTFw5cs8v10Yi53f5WowgOrOWdaB4a8F6
8/K/P+/IOei6ERpvOpKlB6l80dXL72qfG12V0+Mxrj+1s3fK7q4cWZDGTo6+stc9
qumAZoNe1EAWyBpgoEr2nPdesCam3kX59qSdJXnvWuSYHjU0iDPqT1R2aNUjaG68
eC79Gi6rJtyuaG9YASa4kkZ54ag3dBrc4CmIk4Jc8vJiLeKObRu1whzax2wmzXN2
wR79HdvtVympubp7fy0MmfE+Jts9gpSBLaj7WrxmjaqWvMcfhQ05NGsl/NBtmjzh
fUVXFFkhZrDbJkvcmHTPoU9zYh04WLVTERvK9c+HLpwY7ewZjOHuqMMw7lFGKhc8
wAVUctpjRio3rqKiriveJ7la5CRZy1F1E7C4OA5G/dUPA8HY3d0bFq0nIePK8YMW
p7kUBvYHux1XQVE3KRAAvFqBvxKM4E2jxFNYTX1+rThI6CfDGcDu3PRRk5A0QUmr
fKY/9y2YJzlyhTniSxj6cCHCDffLMD3xkMlW1S+89/E9CvZUtl+uMJFqcL6HRrVB
zIoBXeLJ+a5PaXaFlF0n2AdT+WUzwOSUjyXQSaKmdBnj+oR/BvGKzLRc6nO6lHnd
fugNHiZ1ifJMctaOhjnuV0sE3uw8HiQFEArmKwISSnZCkjOqOiIoaZlMVdlfEYss
/w551SSqPYYOCRIaTnSh2Mvvoe+c7kwxZ38fpp/XwXoS4p4BFj2/N270RIC2AbN2
cqIjMzgjmJMZLrnAqVIyOKL4Snpj/l3lKv9hG9rMFxFNwBeM/IJpmylgfjhd9Ady
1QNOt3y+UtepnEKcTyZKX+o3Umg8QHLsrP4sq4NLmYIdgjvhxQxkAM41SSAFEENi
m46gqC2uzxBoJjfDx2Vh3WrSERh0eSOx0TG8mNerO1IrAy5giTrbeoJShnLSPjXN
W/SKuIGhexMAawPaYRlQvbUie6ju1oY4zBdXCDi0FScuFmg+991OpPb77dyij7xv
QIh+TvoM5KadgJJ/dneu5VHKAEzUFPBs3eU52Dx4fnZVbf9fIcBBLfllUBaMlaJg
kN0hQRZeA6NCcD2gqK8EaDIxvTp8pHdDPkfHLL2xI50+TZcOKHUBzmysMd8lVpNI
s6zt39dDrdWGOFae+F2kCSt7Hg8wPlbjtyAoBWIHGSm2YLIQy9E1BuOH6y2rgQck
DZmfDBpptMXq7P3GFejYEbQkFzvqfzm81cim56rZvvazs3J8DUDH5176itepcUbw
C7iZ1lAVzoN/gnTOy55AvPBSPKP5W2LcHjqaDbWZxLMXz2H/zVxs2zsLgFPU4CVT
+MoGw9hzjQQMSJ9NZIKZ4ALA4bxpkf+AdoMq5R/v+HaecMXZyBST47QVmloQ+K0G
oMcD5+uQMfiPskuW0qktZ8AWxDNSO9VSWT+soPl2hXpvTOxf0gKZsEwY0QGbWDMF
t5X0nbEgck2BjhAr/gntOQ436w6gt8Zg+XwhEgkU6FbS022zbAPfmHOQROsi/PQi
HDZJcB/I1qOeT8pt+W1SPNNE21U5QRfF3hhLA22pl3BvwNdBbp3+Zc3ypfraBX4G
Rgcv79FnfIQmyTWCA/8WZk1LVgZcT9yhTcVjO66x6/Vyd27Wn1lcaypQ4Ncr9hWo
/CZOeQRERxHbhe38bt/Mgf+aURDJWJlMsERn9P/VbomyQnB3QDM7zLSDq0Lpoe2h
Vgx3cMazxEl0fcUWnlQ6tT4IWU7OrFcGR31ek9xZWl435XYBITUlE4FcrNMdW6pl
1qgQ8vMm4wkyHy+52aw5AArMxV5+cqWPAKLu7eTdWcgESCVIhdJnNb/74gP0lEVf
phB9vZvhNElS7EneByB+kRxlTXTKB9v34EJjiLU/291oER78eIcA85okes1LlvYW
gTksfM3+h1mo4PPp03GIDE6i2Zr9Sc8ymT93vAvsmLV6B5CBoUiLv3782oIkndXc
ArCkPvkjMzjbFDVdk9W20mJvMsF/Basc5DcfjVUF6YPrOP/2cAtMH3bQGalf8fk6
JUOeydHWS7b9vjFnjTnhtS00kkBba/UJ0FAyUiSpz4NayY1haRFPZcc2/ygcEx49
t0beaHSE7og9hrEfWuD4ekzWly0y8jCKkfUoLZd1Xe/4zBLh+68CWMSo5KPFIo3a
hB2T2NsQ4JvPhf5RsPprcURTJ2PhNHmAyuS9smK1oDO3mvd45Ytk/v8vlstwgfrM
4uCwoKHsUINYo9pqnK01yAXe2aUa3ccqDhc0oKGVl4dudxY4fXhNyGgv3zwPEmdt
GJJF/DEJsbznmjpUNZaNCwWUmZvE9F1q8wc0nXHH1o9yotTFyZPQt+N02H3OEDu5
rEwDWYu+yh79guI0Cg9Zj9wazLcSPT0dmCc44KsCtbhBIR8XZVdTfVIBXaPjaToS
9UfuXsCED7Bo9v9DlAJXM1426BcJ4hI2XTcl9dxazlYuRcB0QVwduMb7nYQOA72E
0/rVakuEig7LONdn8E9rGwZSYNDpj4dJg21HuWBGhKbriKvFEIbG2DM0fUAjtUnN
4d51EdQufgZHFy+/oCpya9fLkQU2A5fYjEVA+rZRnORsSJw0tSWbRELV56DZD67m
cafV2+vCfAULPXH+bWv2/oEN5FUdlx8x240leAsxlZkaNOP29SF4uO8ZQXpHPe2r
Q6ALeYpr+gu+Rpu3uVcXIYSripK0GCKGI560xZCYRETrtNyN2CiIIHoYnM7eYIEC
P/frA/lSIk9q8K+M6JIz2XC08suLgncebz3F6XQ232m6+CdUadgKsML1e7IRAzN1
0VnOJlgYuQjxC4+zGX7/XZEclycuo6J/+ihti37tSF7PQ/jwo2cwH58J0C50Pejy
Hk4e9fl97Y/Gkurfqhp2r5PVmNCRODmhaEM4xeTE9wXd5LGcRLsZjOD6rUJ/BqJJ
F0uRTCtMS0sLIuv8KfPkYJSaJI9q5jKpYY8EChsVDsuBv9WH7McUhPm8K5adJrjZ
W7dOCWoWcGJk/qakew/C00u8CiRcGhB4adnrC0QCvXLQJLUqYlIpqREqzYIq2Uq+
x6UmHzQ+QdII2Uj02cO5PHyUMcovCOys+4KyFd+srxgnMSAuc5d1wfIbuxSKlaiq
35yBZpPGLJa1oPR8uKBcx/mVv1XiC/UP5o8qAO6O48t49z9oM4JGOMGTJElx41Y6
Hoz1kF9iB5dlkqBgMmzF6F32CLlOZIP5QLSOF+vOwD+QuJ1347Jwjtye2VzpCiaC
pO8pAsiDdXymFRyzGwi64UItD/2YoACZjs3KGPp4ycIGE4iR8SWoaYmSddB9ELM3
wXxQZXJWqHYCi+Q6yKpkluJFZmcg7fryEOAjDYLCSjLQCJhdcoJ3fHkuLzpaY4sX
cBDsj74eZVnYSI67Ctkez7scSgOXV6qORXph6tOvU2L9THJqQ+hhJkvQZJUNHCmI
yoVtPctNTHEuTPQSr8ylX+qn/ICwTwG12Eci3l8cONXDNEm6aTa4OfgPcY/G0KxW
gs9Xt8Hnszno4VEfJmA4eWGglRPOMf4sUdVy80Yjr0dcomtnrGjf2s7hwtDYEU6O
6G2MeQE+1NoR8UOQ2gLH8VWnJsov/qyemnUQKqfc3n1GBGG/LIzR1YBXoBYjhnM+
1A4R5omevau058zOKQsBAu90ok6gjtuX4K+YuTn6ZNclpKBkxYb4+1j014bof9hM
PLKk/+xwi9WMpre8ajeg0GRS7PlvRfRsFLlV073KrjXEfLuU8xRv/hOaYPE7VOMJ
YRHGn+XskZCjPM0VHG4eG531maOx5XUZVSEZRrGO1B4d0CwYSnZbj+HmHodFLdCb
ZAiT1TsKHJlwg7Bco3YkRZ/Eao+3OmstHGZQRvyT3mny8TWjFupRoGhmcbYPquus
1jHnP0nF21aKyqWHZlPyVQUhekdUgFIImAWt0ad0EB1iBb0/LEjbIMiEwoTEYqsy
7AprkbReJvAOOJZeJNw+jwoV2FNwtyAhyqloSydDtO9iz/eKIuUVmuSyytO5fJnT
654/Q7VOPMYCT5KCvB2AQoRMyo25IVD7AhdZYGZaJGpld24CFcmJVFolLAUPoE7F
V4NF4zCQuOagNxy4xXWsDcp72N560DRyyT+wWygvoX60SRCjCmPQtZ5WDX0eWl6/
BPspyZYfbSMD83rEywm8159PPvAS41ef+XrbdyAbMqfVP/r9E3jefEjfg0LvVy3e
H/m629FoajvJ+lUlechZNd1MFjscg+4FWK514p4spsP7gB/As2y8dIktvSgMNKC8
q/zTCJx51X8cM+9aaQclGIX4idoCkhm5WXYDdLsi4HNdug66oRn8jkyGd0QNW5GQ
RNtvJAVX7LUb4FICq0/4XMOuWsAOBP3ppptm3eeaNHI2ZHAa0DDgcYbrEHxlm4PL
amumGsqStYbBzzE/8S9EnYEVJpo5Kp0tvjiiQnWBcmDTJR69B64XpeOgHQyWOrNh
WNiPJyu3Fh7hC/oUOAffg6P5awyXaGvajAhBCoqy0XQn13oR/X3Xd/j1JoPlF4Oo
q08cwNrVvVq39odP6s8hWur60M8X9cvaRvxjZtnPdT4eu+b2YtGnCSK2/Tls5YLW
dI3cvSbwsp76oJRD17LaL9Mk8To+lcCe6ZfvYVxZYUqjjpPcmfYVQ6ma5+vC2kki
54kNUQ3sqaepxrWs4fpT2PfmJ7a7unGcbMibFzLWzmXRmFZKUY535KlLo7O6GV7N
g9sMFm0tdMHdSbWmwjCqj0m6r+tTv6Rj5cDoW8MIHHWgXb9NzS88TcMF6WEYIw7f
hJJ2EeoUlAm+MoFhSHagkXtuc4z5flzHQSoxeI2TJKLWem+OBHSv78k5/+1aBuRF
27i+WzjJXqiOM0iDlhflwZn+59gdhsJp4oZXcbPi9Lh/On0chv3xbB8XMzOi6eEd
uqePxAKz4lY5Tg4TeM/I2EUqeJneio6W2ovcoTFGSjoEDVwB/JHRB1ulFisDqDZg
0l+J8hGQJ5ozOC0aNRQEKEc1io2iqXta/0cooewq7BW0y1sMYFJwSFMKnWroQZFZ
aYNf2E2TEHhnCnDkbCvcciKYzVDyKfFNst+aVOWeT7mtnFQC5mWk4NZBcV8jaWOg
XVanA0YuqToZUmjGIoIvOHQCVYBJAt9LjmSElc9xjxVTMQaGewchG79QFsMfA7fx
ikkQOxuSWvAJH3Sin6exJ0++KJmxvQhzhujNL2glcudlBr46GI5GTNXTxQ2lJJlQ
GelxMbp5S/RPK71JUIUIFKVxDl+Rck74OSsYzMbJ2InqjMgX3uaV5bxD3EksWMO5
m2BGdumy/g3+RWoqzTCcwgODOLEhEoIV5kbQPiKZdgDlRy6j4pdHoQoXxDOhMDcA
Zklgmm94B/g6pgV/YuoVK1+PlpW+nSFxJVi/80+0cUC8lGSRLQyPFfs3ugfXX2oP
aRPNbDEvIIyS8y413IjGm4vKxTtCE23FUXl/kf8tOFcOOPyIBaLy/Yr+oQGE3g0x
OY29+/lJGP8YMI9AvoaPTv8kNSmPfO38VvIfDIKarxuasWUbeZPp525ve1NX/vO+
9W2JAlD/KhLwP/gBn5qMFBOAWHDt3wpLXPGZRsiCuWEzQOnLfeo1xU3Id474htT3
p5LuomCoEkk60TrZigiAf+YDjUwrj3tdv6iduIQ5SlBRvheLn1Fd8elxFzYlDP9o
QgSBxdYcvL0eo7KD6tHm6rriGgBl8Is+qCJr/qe2CieB6rVMHU+7Ud9oY06Z0h0J
EmLC83XDHCspIKPKceS5AUGucSkLmiQsij98jLaRBG+3XNFASiBGik2Apkw0fEKJ
E3wp9fjugRZL4FT2nY8oxsm8aWkHsGsif9Jn923dtyNrxxxlDQ+tDaaHMcI/BWLL
QUZI9+TgLNPogdi1ApxvMv3/pggl7Rj5M9SFbQLrDjMp/khI2Tnjqcf5L4w+8bCp
l9rEMLVoPQkBcAwnuYDM90mhWM+1C/YKmXzp4v/FG9Rdjk6Z48tNa2X20AoFEsKO
vy7F0sTx9CA6gUoF+39ERVsAb5Io+Fbk0XqmAwcPa2yUB++NzMRGs5bBci9a+vi5
3elC/pCPE3LxSd7S7NQCZl6EI9HVUsQTf0k9VZ3YNuAAFBuRA1KKtC5OGOuWZEfK
1/tjbfLmfwq4fikOzUowSaW40TmewaGWoqFPfvElMwYlwFmM8mv4zbuNPI2C8Wl4
nSLC/nGNASUmx2uFNMBQuaTZZOQ2dRDUsxDWf7f8lnWpxoaGB92UMXPcGdtzHAKU
pc92eXK+lCBdSWEQiiNyKV8Rks7jLz/7ZUZ8KwvJwZXA9SFWKNqkGKGPPWiHaDq/
jOdggh6P/yxHAvxCa8/ZgbhisDBdlrOvLKld0qoJcxV7FWPDCcE2hFGeIq3gLi4V
Hn6yl6bTxf9TQ5MgAR2y02lhQNYfHUcCv8/xKXRRm4PzW8fDSwZXaJ+1Gs4BAB0l
kZIr/q6pYyzpv3McwQDuvWNfTYWH2N0m+WCVQ3vv2vQUhDgvbPk92i04xwuZ+BMv
jVMOPPT+GzqBIu02X9lb+Z3xw8vuNNY6PilaUL+DGQyFW3SBjZrc4w3YuQCfX1cm
aFaS5MTSL38WfHtC1HQmrNzgE/uw3iieWkQ7UNyT4og/VjqedY3isiO3irUrEsyS
9QIXRCj96qS3KtyZ1Ba8LrOV9Nb48NtFSdiINuuW/aWO8DvQk4Bfk8aeF8S6kjwm
0zbWD8nxFshkpsx1YBUXMII3h/PjTh8WdzOicmwbl/f6NRjKkyu2yv9tLVMqlGvY
FpyhgMj/BBUddBBB6f/d/LPhnfETpWQw2XRNsmJDD0Go14JsXJo5BhtVZXW++kHn
WnF7AV/hp+KQs1V3i4zcqbVoTADubzBgYk41K4KNuqzDKtzBVmyTEApUAL6W8Erf
/L5bo1YQtND7ip6cuxgowZvWHEDLEZ6gm86c7AkkGF6LnI2sNYNmaWa+iIYvwq2u
2KqVej4bgzfmRQ1BZqWwVFBY1FHUSARlMIRAul1ZZEiVFhX3G+5A93cwo31esTVN
0ryr+Ja0t1tsvShgpi3tQgBjgVfoetKF1rEq/GkHIGoSw3uhSkJRbzez4SdG+hD5
xvrzTkVYvVy/VVyw3YB4zExw697a4m+h9E2AottUHrY5Lk8C4dtMMvlczPPGjj3T
8Bp2a6MMgXvZI97Om7mvs1evMzaryAJwUx7BOuIaI60Tu8uhFHDBTCrEFvjHrmse
i7KZGtL09XtqoBU/mn2uY3F6S7dsBSSLrLUARgn7vpODKaZHKzw+//33Y7JqdOe7
nY0f7VywhkJaYS37IwBWv9af0Z54NvpAo+yWDJOFsxav3mDVtpsON+UA8yMskYPT
Dyhqet9DAf9xrtrTM0w/hh92AjD3RfUwGIFfobNL5GhuSBSRGR60VShyiKQJpT1p
10ZEPPawGX5i+FKTbscNbzyaIBGr6Mv19MjiDo4+DgL6knCsd5pnjZpYGtE2L9U0
ipcJxrZAgYCirKCzSEFHL+lPAY7U+JyDRIXRrMDRlLubS9RaI0yCK3Gdtt8/G+fV
WCmP0crpDXRSiFsXUleIcA/8rY/B4czBXK3CpBYCw7IPE00Ta1Hvz9bjmIYcS7KM
/kfeuNnkR3Ep+m/G0xwGJxEKfUJzst2YAfI8It3ftIKyR0kf/flYHmKPkbjiODJO
kepDXs+fmkmDMB5zfYtpJyUyl8n/w1fVVQjpOphjZO8CKHzrycpanWJdH/k8/LMm
gSTQpsxT579nr8avfW2bF2uc+/OMnIYUfQxInwB/uMydcbWUOjBOvP/4sOpfZE96
poxHt46vBDmQPdin82V2MW9S2LkeiBeLrAN+D5HGaOCYWOJHYMS6j72f/Do0I/SR
AUdY9OJmJT9Bgc1HVQuBAhmssAjusv+ElmAInQumGnaBBuYVSiOaKO4s5r57PBCm
lAEHCHvZWuZ7w7WM8S0OCUBvjB9QXlrF/ftBRcXYpSztHyHTmqMaSnfRvGtuKdOc
k2yslJUdsmrtb1j7hND9jGVQoWNeZXo2NcAlDu8IjyHLODWnsNWxG52HTx7TJMGm
tDKxwA7j9nZCD2LQ8mLd4ddFv2lXqDwVocKdfU8KXjx/51ONfdpYKrKXBwohcikh
jP5itoklg6FffYixwbE0l3nBEuOsqCxM1fJIYioLNNUG769LnOxHB2hhGZbzDcip
Oi3+OQjQX8Bh0WhZEk1L2GvcLlbGsQU3wyKhbcD/Ts8f/6zR+HISw0OUFdwRunyt
XLPcOd27MXk12yxp5O9gxCpYr1s7W1DfX6U/l6sC7uC2tya0bWqTdOGE5FQgjzaR
AIuh6RJmZY7eHyy5nSaeuaP8/GQj2N8ZEgmcrslmAUwitHdbClbJeEPqXZXnHLUq
h7DlVvI04WKXP9w3e5nmKWQmVEhqq9MKH2zHabLcvyMNPnmdWyJnH8s0HyPTbN+e
FhXK8nyehBNMJYlkEe0R81gpI6EB4GF7Z9YgMBn1RCaQM2jGPCWxsi16FFg2RjL9
MTUNusgjvHKfK1UK1vumVeb9ZySW6jTiTO5JwHlWtha8pZiEfsLy/ijjrLqOV3lu
C82GXLjjRmm/99lFcEldal+A1fLPoPpXL4T5uRlAZPKmhA6MjXATY69PXUR38ZJT
zwY+QW41c+jBPUjjPtAFr8CphcfE+hg3HazgmHLzWyPqqSS+5GtK2Tz0BjReTUnE
+D6IEBp1M2w/qZIFy/bgXo6j3blFHMDhuR06ar+QOYa6LD1KBARAzIUyHVkPt/4M
sdtWe7u5L+GBe5A92V8Q2BYDy4j8NLg4t+MwEBWdE0i3O0uX1SbQtBVZCLafEFrH
so4o0dKwW0W94m1facZMi/OlVzq0/6hwindCTZUbr9ImaFNMwpe8CZ+zfwe4Wr90
ff5/BfAY6KRPQEHlgGDaHjuZLbZph+nFL7CtwrpKpW6DmIu2CG1zPugWdQAWX3l+
IQl8tAjn8qLo+4IfHrjRiRoDN73AL27FToLorhgdhv+fBdWLE9MiUj+118izhpcW
zvd+VNSBqafSvlkXrtjhO+jL7z/97uevaFYcdfXBbVdGIAEqz0ltk9WOQyA016sa
VC8DpVpWoWBVvqUbBAU7FLfdZ+Y4ycSRwVTBCJW+IeQFncSHpuCuOHdoWgw9i4Y7
p5EXnusJReiaIr0+M80XiNJ/DstT5dUqfvniuc+RbMmWjI/RvUfQTppjvDTYXeDw
pRCa1FehN5HpNwvnk3xd9KPjB7fHXgf8tqu6ZVuPgvCrGmlxaZwHdua+3Tx7APZB
kxQgH8yc7z6e5S6tQ9JAzUda8J7y6FV2gPJc3Awt+I/Ibe1jaQVOUKkdOKdjSOSG
9CLfvR362EN6UQLEV1rQdnzchpRT/IWUpVAR8Ri0zEaUthqySw1s22idaW9ydBoq
8kMpjQwOO7yDhzisn/4xqWMt5nrtMJ5Hf/H8H/IzTeJRMh2L2fgoXkhTZHOmeIaA
zbRxMDpZmTP0GRFKdjJ0YOKYODLl/6Mi3B63nju/ms44ceeHtljjvkWTyVU3cULt
6KWg+9TSBN/dcfrdezqXG+NTJL4U6Up/lEotyauYG0CJKLJ6FErU/LX5q1jpF/6m
v47+U+HfoOXkjQ9ra6gcg0wbK2T2oB+zG8yCg8ojGivbalxhVQ0fIHg6dYLxfKAJ
S2rpn86/NvmkW4MQnTW2neGdMP4Ppv6tTf7ltXBvlMnn39rgO12R+xXjeK3quB9A
RPNcMHB4pi4acE3/D/LCRKueo2QbrniAjSzbRdYK4oJRcbWhpazhXxdPGiQ7jJD9
f/eEmVEdGj+YdCA7t1IjPM5j7xmDBp0mhwjxBGIenP+e5EToPgB94ouou6N7KBN5
IL9XISZSeH0PYuKeN3vkiG1ZBH2jQYLy86B1XWrrySEbyUh48qeSzUwbqAXa9K4H
X3NVkEA4AtSn5u2xGj1dC9RGx/pNC1ezWHQ/6gPOEgmkq+DDuQSn9krwFZGtuUWx
/rGLmyLe078o5hzpXpStEV805V8qJ7z3OPFFtzmYoljQF//PUJxAIUPCFDOotfn6
LH+gT/aZLaK5lJwJECLh78GzfUZNrVV+CkL5URA3zlNUrpdfFRS98reblX7PvJMM
yhszUWv+CU4gg48rVDhXpcAgw4qgIJEHlyUxScAKUvgN7f8UDetm6o0C3nZETsT/
NXVpZsajWICGwesAbZsEA8clssJe7Ym8GKb1cSj9uqtAEe2lpj1MLC//tBQ1lMJP
j48yu6MpOZkUe2/0DQy6nL0VpQR108hlAAtKEdNp3Aek2YT8T/0+UuAKN4EbEp9k
Dutkqsd1eSQepqI2RJh3bKnymktf+S+m5/f5KCltyI0P3Pt68wd3lt04IqVlgl5b
ajgjKYq05kf0czmcEJDawN7TQPliB3alS+rVsG4w/abaJLkbumjrg1rsXjKz7XZ4
qfW6h3yPFVR2epfZpHnmv0qYN3IzOLmp5Mro4cP1BWwHM9f8PjkAKuLNVoGHmjXb
ViX/G63qW0Ksk5F+vNg+o73KL6gGz3GbtXyfviv0Pf3ueBufuJZEWNEP4UpDYWjJ
kji6+KuI8MYGDY3mqFSjWDia0OZ3j5+9UfcjFfnfrIYln3tnQdKt9KdWMurA0fqb
+ZEe+MLCS94Cbuj4Q6+iZRo817j77hxugBAKtZ8BFmk1Lj6ZLhezYxW30H3sJlIq
+PyNQrOetVJ/DGSSiwvCZqqbVQ1JRD47eN1NNzpnR3mWeVYBVSkDGWnnOX0WITzz
Y6wMNKBOPXNysh1lzXadnv9tkVVVSJBTaM/Lz4unSB9H4Ga6yIo+WKh9uMuNnn4S
+9e2hBPlxEP/8TokInPVN2X5vmrFPNA0KrKs+vcV8h4zNJTGuvVzZkRwi1VEfKBF
6UDDWq8HNn6D/F3lqGZY9EtxTvIWIgCj7HEkNu8GJGD95K1Jox1UUazLvpJDIyss
Fx+3Y3QQSwM/OXMr43QXmPNqzR4uBrOFeBpCU975bDrpXtEeI15gLyesm695oBLZ
9Fk4S55E+INadRH9hOI1/qAmqr9vwO4VZ9cXCml1UBy7q3XE5DoywTbhb91Mjw1Y
J3hxmsNMaYQVieOXShcghEF1OJHg/cPxIkfGy20ksv/JN+SHxTqOZ41NvITJdQQG
Txe6PJBRSXWHlmVlBT0ghlQaKu6TLH5ps3vt9Cm0P17z6CCuE/x+FCZMkWIAJVK+
DwOQ5RLbNJtGgrdOQSesbOmdgKNOYMb3MZde5b2XOTzBsMRev6Of6MDjBTV7/J/Z
pdy14N0CN8Zc2CuzO00ck7LQLlS6q7mVHu7Gk878GMjmSFeCUHk0uTH9pMKlskag
M5y93uDJRUY80I8S3x+MrguzTa5uA47msi+GR7Mg2YBO+eBieIu/BP39JE8rO4JC
w3+oyLeb9nf/9tH9dNSQ5hGUTNllsywlSR555p8ID19QAztrhzOj8ze0aQO98d93
87bDU1+X3wQwpab6oacfVTEHY1bPlqKkambVSjK0tmhG4q0d3y4S1PQal+uu6CoA
LHDWaT0XCdsYqhswQwOtRRdueP+Yv4+nDeXx2+RkTjSlUNcn6Qq1bnfot04Lkjrp
9oMGHK0ccRJBjUNukV7Syg4kTeFHi/mnVO6n+KzVwuc1t66GX1xuw7h/eLrnzadg
TzxHlUz5D7a1ZFc03cPI1prRAuWIBtsEz9FG4WLncqZgvzcaChjrq4lpukaYVb0N
i9zOnPd633BpnARTUCFLYyMz5I/O4uy32YStPVHzAS5TWX4OEONzPslj0u9m4D0C
fEjU5eSDv4m1acI5FXAY9MJxsD6G1vsQCYRmhPgSUnLjgOfIUQloeeaB/n5p1yVP
nDEOM6G2a1vMLMyIhvIxgcBmYHRRvp5fv6kJoiZ05xfkNqWmm2lWCuHn59Jc5ywA
hAQkJgxX05Ut25AeOqq/Zj/UsPyJoi4EaqOaTbrg+HkcuE3h+hYvJDqKqsXQ5/r8
TsL2dHFryE6a4oMSr/Ks4RGSZQo9GjS3fpdq8nFUvZX1qtMRmce/fyjc896Bs19w
Z06Dorj10UD1+W/A5cm3YvF30khNcf+t8fLSz7GOf/gwJDtVzxoIP3wIs6wR0Jkr
DM6D/vVPewdDxpX04GH/rKUvaznwi4B2DicWHQj1LK1T0G4azJcIC/P2AOev/Li0
r61dY/Z9FDOPK4dRprG0M8EmQaDNQ9vuklYHtBC8V+nKP3rCWxXOMle9hWjbi6RG
VqD+m9GaQuzuSuM1hfWm8xYhFpt/RIX/pYdYUKqvKgz+7s6o85A98tKYEaoBk7EC
BWMbHHEMy8fRZleJ8O7ScTSa3yMEomVAsOjC7tZokFCCg8gr3bDDbogydD4aOCYS
VmUrRvteIgpci1TYBkc8rZBSXexf/KTIzPD4wEQRjbyVhTPfSZnPGSK5GdhLhp0w
gq+QScwirrvaUuvScjpt+dJ7M7VW0OXMIVYnL27atIcHVljfibvyaL/Y9UeOfBLp
MwMsO2Fifp/C7RDOGjFqS5V8QgsrYFmVI7pdsfpUkt399Z5WE+GJsxEM/X2emJ+l
q1DL1U80lZB6pyiCtDitldNXsdhHgz3gJofNI2Gf+3TQlno5GtpcTmWAVeFJcZ8q
dQOic0F9XnprW8Wmw5pJFAkDjbRBsuWAmqEAB72rjTPc8x43IlC5G9Q9RIj1hARF
rS7by79vu3PKCVDNpgbeuWZWSsvjd9KwPmjQXxmgsp+2LU7K70qPqJG3JyTg9EQI
/x9lUltWF3Ll3aY8H2I4w6HedWmjl2eyj/rkQdFrFjbpKpjnkgXE37eX+EGecAhW
nQVmhRZSkc+OC1336wn4lFL72SAgqC7c+lxb/RjqJyx7MhCadDrfbRXXcOdYhkAT
8rTr8dAGwPMatdhEete0oyQtjs3tQwjP5IYpjjjhlgY8+gInNB9H1sUXE668VxbS
eALEGYXhdK+vyIVuZqcXYcHhmZkZS7XpJUKxuyYhwZCCLARjidp77m4F4JrDiSxO
VBQPN7KlU8qFcK7d6QgF9agnJ2ldUkAAIv/Po++2GgpuG/mgvRLMM59WgXOp3yno
XzXhk/31lpAMIV/HcmI1Xf4JYuknrbhjOvz9HGapDUqfkzaI9XIRvjkuVsn/8+SJ
4oO6LRxN+8u1NKLWWgEOf6de35+ckkML+dJpF7RORS3pJg62N9rJmZ8zZm2TCZsx
1D1EBvte4z5vcSYrvql+dgz6gjeQY2s5tKIK07TPYXEOr8Jh0qsvWMl2rM8B82G3
pkDWiPL74PVanyJIeCSEwxbfldUrt3qCRNJO4AmRDnPGHOLYKxn938CZ//TzQ+9L
R3Zy7rF8DM3whbniF1BkwDqFm5LPNlNLDhekZsLK0bU9FwlECdp2TLAWTvHkeRLL
/AuXSrrJcKLwqVlb9bRG5i6Wq3/Ubt4xNyNNLRg6DFPZqhw/LuwFvYyDBxobPJrc
55qAS1kpzNSH4o6C118awdMUwQ5YMQA46aUsxQGbHx+rm3IDMHNFkJPLzP2vtKMo
EEHOB3Gd+2/+lGnUgTLMqx5GpgcNOCLGe0UVv5CkLXnwP6C6ZxyEjeNRDvNerMYY
AO7WEcop7ZcNyxhfhuNC2GlMo7rjNRjc6xVEaSBdp+7e2IlwmUoOmGqZLB2c7Rb3
zs/MvhfY50hDE3mvAVphDECKaZI8oc4GgUzuFzggaVYyC/kc1Jggkanxh/+TZyLy
aHM0cBU5nfA6Z0SPWyCA70EUQ+9uEKKFenYDu6a7+oXKEod/BjAcElKFH8HmettO
NdP1E0DdMqdCBNFxWW28gU0KE9bKPgjF0Uj9LD0OL+SNyt8ZAE+5+Hyy+c6k5bEu
uGL6YK4cLIKHOHiV7sCHwNl3LUFTYQmyg57alCMJAfcSFosKE7nB0cF9eBRBohNL
Z8SKgV+9kh+TujbzgsFzcwt1JKKnhW+rg4z6o0vLbpg4vnDe7k4JH9MS411p3GuP
pCOkeBj3f26OCfW5tDtYIGfMvwSnukith88HWaYWYDetQr6xYxFFO8LmQjE7lGak
IbW08sBINHEHbVbZbC7I/zPA0ERVxnwW6vFZOyWav0hYoctQqwQ+DAKK0vuqFdhS
wXXZPno61AArGvqvishgeMqOL6vU8hIt9SDpKHEDF/hBdq6sVQLaTedm6B76bRFo
JNhJLJA1IDo9T2qbKEZCtFMAj28T/7dYI226qdyvDPYKZdrGSQhr657vDOEUL51v
fnkjIHXYGLXUAmCSmiwtkXUBi+CVvAb6xtVm/AWaz097kUqfjAseAH9+M0vZ4dqK
K5yZ4xFvOFdAQ7ap1ZGMl6DEC9asnyKnrh07li4Ot+ai/Q5DFbSuuOlu357AgxCe
7s3fksEL5wbB8YKeYmxcpwsHW8s5AOVNJc6g0zQRw6o7e0CattR3ejoMYwqquyYK
QtCI4BYE9Dpzc0PEPqLc3pFVpxLJ9zOs8gQeRAzr0Q7Rw+slnwXRA4u29Ypzwwpe
MlG26fCruk/1ORF3OnVEzADuNY++wcemsw7/NyBkG+3r6Wu17HAKjruC4wrPYeF0
qAKOz0l7pmf6HT/5o316rGX8ATdtiEd563K/NelOd8tTwLrASwDo6HIN8Sh9bPLB
wEl6DmRietbowNnsl9n7z1wqrXskDDv3qDzTpKK3CBSEf9Bg8p3ratI0CqHNsZQd
v7Y6IV+AnTj9SEPph7UF1cqYzJEl46vhabwuWubon7S8MRkpbVg4dNEO2/7wDPYH
bVDIIJujL+WCyVWBynVpOZ3QT+ilOEJgJqga9qjasNht6LDe9Hx6oRr3KCm8nJdP
XhDK4W59k6ZnmKgqhJ16v/rv4PAwi6IWSCbmqLORQvXPhDTCpByysWzPKSlBxAPM
4lZEdXd9G3jkdI9d8BXjoEY1PCFAU4vD7hZjtjZDZbpvspzZ9GgdwCagaKJvIdBV
QCLyoCQEKlAiAOwUJPSxV3ix1gMdlasFNECmocM/4MNKxJ7AgJBcynZ0qxDD5pbi
xmUepIH2ibQ6q18bVlWP1+RDe8fmx6EPlhW6ZeNp5yqQjrsBFYB+o44JRKWyRed/
vEKAHm0MyvwMAOyKQqwWUYMnc+FbWWRh0qSt9nGg22VN9z0k145s1fQP2PN0U1it
0wWc3JzvcfFu82p/OS8vBkjxDot6LgI55kwWBQlLfT2SVvtP3zsseDZoA7fWg95W
gPL6ThtNnHV/Cif9Lk/WPzHW4Fa5u5FylCeRpAC5YfQP6RlXIxCsQu/cFeSMiuBI
53Vf6lNgC6GQnyJ87GtLnw/kQn9yMN3yU5WpJ9lxOpTHQG9xPDx2gehc1dlhMxTV
cdFMN6nzM7aimfSKpVVczzX5S0Gv1SGTgsv09V52r2GOCpoZhc0mVaUIPTDlMh03
8OiYRBI71AZjISI/zZuoCD+rgtqx+CjsuyBycJ7yn2tGNaiZNxlC4hkPsIdBe7Jp
vBJJoZeZsqooq8zMUKpePd7yai9BdvYlzPm1QWmLDr2Ir2FJpHNARlW/IB/jrx3P
b4nPgzsns1AHM0j2MkwNPwQvszKxdlNtOZCqcjXAKrDFzXMryYN44aVRXncC+z5D
URQoEWD7tY6ONmrEZ06vB8nH6EIPdnEfxzav+Lhv8pNkB0+3OScYY9p/gKNJF4gu
+TGXwevzNsquDNqUZpfoJnMPGpuex6T4ehfEpVp+4fbkrheb1Uh9NokBRzd2RFip
jYCu8Id+FXFxGvcR4A3IhNa4BZwo/JYoYJ/FT8ji6EQrRY54KxTRgScBQn/GxzCM
9DQX3MFOiCj9gfs16vOk9reglgYFXGA+L29gq8I5ZATTCLIHqGxNQFTmbCQDDIOt
w1t2zMOIutenWluCjjkrUcjcYT4A6YUgWw7j+QRfFHmIqHQCjE1a3gUAd/PyPERM
KQf/pVxHmTPX0P/OUJYJEDJAq1Sgw4nGefOYVErHKGxheGpb8SSAoU9jkflKF7fV
K+2F2LiFq4ByeQSWEzNgiMH7n/Vs5NazyZhOA5y3crjwPSTxL9EvVisEAIE14sLO
Z8NCffbZX6POOheF3yDWsK5kDGrdWom3EAcacHSR+QVVpXMcv2JO34/T2/OT5dU5
csFzKtgGbPx4V1gDiiTpgOsnAAE+R6LX/usHzANWjdv3+Dlk0WtuUcmcHO6t451J
hkhEE8ddQzdp0ipX/Wd63KVaQjXgSZuOu0SMcGuK1xAW8bhBCqZdp/fDY4p/OJmw
ZZnLOT0xhv9XMZYFnaa1Sm8iNnW9MGso4Zt4CvAzhibMSI/NSgf4JuiuZUBR+tOK
XG9xEWAYNKFeA8/8uqIDH2MwU+4mDsPXO3kIREXSb/ontm1ss/mQ9cYxR4Px6Lhl
lo7D8B7BiWMZghQGt/Q9B47qFkJcElA8ZLWJ+CN/ifduhFcvaKfyNTFo44vpJfW3
ughkwq11jaLtE8xul5TWwNPT9ds0IKZJg8KpX/i4ICsIZ47AZgUgU9MAPOWyPK/3
rXwjRbNokRmuloXRFKMeevdnbaqIVMHwcSxItdnXokYZV0UlNY3bRHDTd1StL6ud
M56slq4KT+r9wSjQo0738UTlyJ2y9sXARzYvOxQmNlSOvLvOSoM50liyxsJC4/sr
7/As5ElE6um+m+w1kuXt01FRgyfBPaqqSW4tOnN+dWPlfmdVQsdjcTdJsEi2AZ5F
ZLoY9Cdn/EOsvcZIX8RinhnSs34MlJkWqkKL6qWk/wyub8Q3LJsVa8832vyQh8L8
U2DsAEVWFXqLu7FARpEnPHN8nXFl3vtRQAWxUg/sFfmbL49ETKBK19kUj/C1GklY
c0XEYitfjij5KFeGKZIxjCRxZDgH4uDtw4ImFbGysOWI2BYiJqYouG5pYIHpge4U
Mk4S9MfxdEwneuG0SpZ1kMc+5/kIu2/fm1UtT0Rbt+FXrKJQ6z+NX/fEZLdZNYBE
axiX42817b//n980d03JL1N/BCiZ+rpMlS+QDENanpOpZowJPQDB0G9QQX7+iFDx
2/ya64RijY4ITr5FFKJNwzyzYmQvWyGSDuWB146e/9ejco1yLPwpsqlPcqHFnHBA
VVPS2aCSfndkGfOwIXu0ColGaXJbSfGz0hBm/ougQWQ3SqtiFU1vpp9QxNG2YVna
UfG1AVGGIFcngeqiSL3Tf7d3XTWcovz1Wqf4gGoKHQaDJZPJK5E9QFmKwEjDCF13
k8UKLTDAYAPSOIcCA0PtIXohzrx9owMoNh5+t1hnNN2mqmWWIkPMp0peUk2xRQbs
UQ0IPtOnjmecKI8l5X+eBHU1+m1LG243HiTIA0n7kal0TAlZOcI9jNfbQkATQlTl
rzlzET43q2TeEDsnCWtlZh9BN3/9BC1p6vILLxV3WpwgQW0NcCmGGV6VVJqGTFXo
We7jYqhXiRN7v/BjUnTr9BeRlZ+PwmMmmSZdXehq3x41R5MOlJ+LDrH67w40CLxQ
srA0NzmLXXyfn0C08/COZMYNroc+kFd6IFDf6TWuop4LrKDJzqq2uNA0zxd9nwUi
aG9ZKfAMSUmpbuTV404D2AXwsSHQ6d/P863O49Oc3An/OqjYdWW73XBEW1NgAfGd
H6VTPlYs0E8k/Oa6nTLr+3fYIe3IXUEkjAhwgl1JZWqkAmGinCaCx+3hv0YTKyqq
jWF2WmQmv7y5N8fjRNbnTd04LjyG5gAAkA9k1QDHTfjl/iTn5+6Pv8bQIg1rsP10
yVKnKNxKor2ZqOPJ9dWh5EX0xRKTi52B4m+iMACbd078e+E6B0KTRmHNbsi9QgCs
5fdDwmluk0+FFImkmSTTnkTm/qgIs+5WSGrZRklnmpO6UDmP1EOOcG10RRieHoS3
NDG0NrA4iUMDKsI31+cjqjTr9rUG2URzYlWHin6cymLxsu9daSqyypjW9X7D/u9V
Ii6nAI9bOd4FrhmlVGDH4ANfZsjTI23+imxze7Tk1sbHrdz0iMe8CWz8ZM/OYfcI
7ZnyT3rtfU4EtLBwPN4hCnkcH/jrILiV0/Olb8odywD9NFb5hTyxv+y8oHWB29GR
9+nH8r7/qEmQnRqLbQ5hBprG1godswzKK9/IXy9i0QRuGgMRX+vcB/bM292HFBOk
Qs+wKde4d0CuvtBU9Am8wNDGbF1N0SPPBngGhztXg95vj9/XgQtw1v3mYWRrap1B
dT6jrVYeyWSzxx1ZaqobG483azK+8RWpwEZXkx1RCld63bC1oli3WMbYnbK/sGIL
LNdU2bGcNVAV6pO4F9/RBHO0ToMHUGJVhMmXb/shNkHzoIibcmQ4vpQbtf1aGWXt
gzYNPuQEp6Hfc6NQoyLEA61JVrDB2rKAKdegX2/MSDt3aSuWyBBtJCxYOWl6Lx1r
F3QOAfYRJljciZt6+jRtueUs/Ikyi9r/CoxZhsMskLzpkn5SkpRJf0PIY9favdv7
2MHZoHjZ006D5Ic9CfC3TButmg4f0v6AVuv5PqMv3G+oWcdN1DO4jkOQGi02YK2i
Vv7PJ7x9wA9JHF3QP+8Km/m+lO4xCfg/HM1DJsZrs9VFrjrHPBudLZ9qNr35GeG3
brLNxVFbqz32+WWDajCNNP174YeHBK9MVKW85LlQcisb9LU7DXsReYChm4MmJTn8
0Lh1ZiXbUyAhdGB/UG1EVPthX4Y8fQ/FZgwh4uSjBI/dv0K+tzOu//TSumxabcT8
ZA/m/EiS9YDstcF5K7H0OLZYDS6WypF/OARWqFiVjVnTYebiKNNrvsq1eqVNOl6N
EP7QVNOsH/4biEGVFn0KMlcBxSF2wwmQuZ6uAYPMRERgIYGm6Fa7fQ19JSpIIeH2
j6rC8OYHEjFi1DIScyq/W179WGt6W90Nr70ID4AA+FbnmVxawF+0iTXVmLfkJsDy
VTpSKD9J/8dfh6FtLG45+iXxOIXiarziF+eADMcgTLPPpVmuP3UPhnVD4dBSHc8l
9t5su8E5RNf3yxZrkpAbINxHsl3IWz4qskK6Tdx2giq109ssO7sHu7lWPcrYmyiW
XUhKcVoDIqCrQmu60I8qU7qsWrJ+FR05admHJDzWrc5D/wIHQTn83QJYdEQahPrv
o6Q9JHrvD3xd2VksVYka+xS9TGF764bU0XjXrx0p6Q/fqtYrdVRmh0YHgM+vNIao
6TQ5wdg0f2nxpFWd2XWbWMxZp1pEjGbRqnAKCQuQ7yOsjOEgloOsszTAv/3Ubs8y
AGluoaRB0NIDoOSg4Mmkax6eLR1mNY2o5kbXInR/exGn5lnZVmnyZMR1pQf462eY
MIjY+Guao/1HVoEp4g9zZN+nKoYLA1aR7T4Dmzs1jdB5FieJUC3Jk9nJdg5hUNNL
i/70NgdDIoixBvX5sC1t8yMS77uYmvYRB/SCYRVM81b9g276qkOoD1b4mbKYzI84
cU68iGAKcK0pzBX74gzOvoWrG2UUY2TXptURqsC3mtnrwuZQ/oG4CrtJkK4WnY6a
X8V7ERy0fbHa6nD+w+xxOQUM2JSOfOuLDKgDwTynqp0MaMZmXbAbanlnEcQtcIfC
QRCuwCxGlEKZPDdaksFuHuGwmNswADEtqcFmuSSm/wvSkUGVb+oHowywJ94WanOj
hZZ1HbVcZ9qDyonDPlTFfP2Af2eQlmbj2yQB7Jk34x2A1vIFdyCGiYldqStAz7VM
I6XXBVdUFqstfdzEolcxfexhqavygQ3RTzeEmonFACN/gAlazEq3EaGf5Gv0fFq9
nJ69O07VWHQaXfYSn1JawZLS3TXbQe0VsiWbDIiu2tfaEdp6dhuXSAhhQHoYFVDh
4hH5WdH4/fLZ0fmxUuDU1KUvVHDbD2052p75/0GIAQo4ftPjodlpkz/rDOWN+rNm
HtfJiA4c1jfamUS1ON9ZxXNouJtc/6aIeHz9Je8zLN1m/dCvtI0zYgDQ4i7gz/GJ
nWL2y38WUTKie9Wnex6M+aj/nF3gVcPKlU+XAbZ7hDQ/KKOHXch5D2oBJI/cb2JD
QydypiVd7OSESHXMa2JZQSE2p/7a60usffULwKFI3yVji9ulTgnasBx7q5vaUD11
cpDvtWVjR8IHYNc1xw6VBB4ZpdSH9gaVyUVTldNYaJFENx7aMvFJE9oJR7v622b/
QHoH1ogg78JQwyQamocwSKz7+s0qqMjZ2THe7gMbPSqUuMjCC1Q/1xlS2jS5rwHx
/KlccSbQ1EEHu7AwLtODZnofaxdG7g4hXwhvA1ulFNHMUC5kN4zml9W/pQWBJYcU
lfQ9WpqoPtZYsCxaSdMjSLwh5/5/1wQE0QdeBpZhGCBku6MR9DX/kCajkSS2Etxb
DjEdMDp9P8sgKO9OwLFaUbEI4NCpCLTEgNE/lDWwVvu0P+Z8REs+i5518nXloNKR
unwo6kmQDHB7G1lHYTl5cpHgYzD9ljMHRgmlNaGbHH20SCXF17/k1QCbB1uQbyrT
7ehEqCQDIR3LcSuy2xqRyuszuvuR63TXy27QS5t2tM5ZIlz1yUxti56Os7oVhqBk
TLTZjQ39pXdcxQGb+z4kKBPC0SeniTTIuAUIyWY40AFZOZOZJPRC92RrpnTXCxNm
S4hvbnkl2gyrjXQc/QurVOHxF3yLvH38uoAWoauX1oKCguRNCLNNgh30ltDXMeVa
TNoPFfymeW3Xu1pH2inOhDBS1mBfsW47CwCPS+mEDi5AjSAXMkZI2oCtZMg9spy/
8ZjXjIh9RJ5gg8yb1Nv+jyX7PrG4F7lP+bpqUQqjos0N53pw8i6xj8kyycWNMCFp
hiK27Cz6Eb+gf8XCHz4dpdYhbhIeHeorBeBJS2K/xoJ7LmFyESDRrWOHjTSGqpze
ZIYhvTdUKRLn/xI6NJ5TMp9Vvnvi8elAVFIoSx55wANDyIXS49C1cBfXzSsC7oQC
9Vu9R/8EzSP79NqZX2d0mXhW8LMdYPcrNXN1M9kh4uA0qI52xAK1FRgiKI7dzs8/
6ZL43Pq4p8B3LdL1fP6Uo/p9IqlmpWAKIt5jzApEb2+mdOnj9fOwh+vhMnyM9pyU
Bb9LTMFEXT8cNzJElcppT/t8pKObNoZfjeWzROZ31CFJaIfp9dckkuIteHetYcd/
zKTAGiciORTIz9dVP3IcPyo/GUu6BI7Hh8A83Tv4hTkbg34hJdOL6FT7KU6og4Vd
9gf7h+52afkHTqVqPnAlL58l9QnVGxx2RxI0XRSb4uXZ0Q8VKO9wtZaNNkKBVi60
DuGJVNQ9HQIahSMdOcifiWxS2GUdHIJNVQkI80YvD5OKv92zOn+lDEo6+Pc0QheO
rE1aBXNE5w2Pn2zM4wcCUS5Oy6/ZrguBgCuGv7pcVf9/12zK/8rPP93WL1wJET6Q
14PzTxCFLVZ086wpPl6pZJgmqgdilcV964jxIy/P/nEzYv1Vx1paZocL8VjjOWl3
eBxcgT9ElDIy64MZdcdjqrBG70h0o94mwPJUjpkIWiS/yO/jsuIuwbVHzNPWukxG
enngBPX+//gSgJpCb+fSrsmH1ynWH8cw7gq4T6LNDw74RcPkJ+JuIpHHUp0uNSCv
VP0NnVaYQzmXwRnM66r4H+uP8JBMdHW5/TKAcW9CwaTYqjxANLNT3/ORLD0lmYMG
WhafnNopWQ4672LM31Ug7IYeC58etAd+VrJ4Qd+ZqNCIWe0ZqNNSPq1E7JE/2pRa
ahgUoosrNVEw7uLY8S7Pi6EYE9WU9ROdtvTmOZtMfQZW0J7tyXs35aIo4zz4SFn5
9+nZ2fACFrQCR6cJ0cOIVhUDqI1uO0OGbBzMXF2+MyaJtnTa73hpJZysSdL5eyFL
SwZvOTCzOHiyG0NHxJv2j+KqwT8/dce9OpOC9Pui3z+cNegmIAIHF7T819acA9Ay
CmUm74Z47PBFpHTSR584fwzgNPiAm8IDi7MveixHUjqPMMkjLtTOKag2Cc8glShQ
vsK8hbttF8eIdCE81k5q1gbFCKYP3+UWSUWhW0o7PLuOksl2QpbxPziW7QroZEm5
ezP26VedCQX2un2vxfXfbMllHdnzuuX07EDrMzqEM1zpzumUL5hnSA8PuJQTXMOn
pM51CELh98uNICgzzgw+zL4U+od2wTPhaUk3+Vz8WuLPmZtJOsMyPqwNlouweE84
DQceLn041Pr8y3lBrb+vOmOMErHAt/pAsBYaZyghNeHQy9KtK8KwNtXczgHZ1tUt
vPgo+McDvutp+vHR/PSCLj8frKvplhZcuvHGtGsnC+dNNV4c/eY2+j7/s4fHFWZi
k8HjFfae8JFjQxCWKuBjltElZHMmjxNHxSmr1EK5nnOCbRXEDAHS830IdrNkkyE7
7OCBnmICWTQHaREwHWBrsDuFqnMIauT8KxkCOa9EDgWkGWqlzuxBr288syVRb1Zz
JVneN4ehzfj+ADtvoauFHVJ81jVi+UNyGxCFYCKk637SnSBFVk8F6RI/xtYWvDlr
flkn59vjfrubvS35PGa/lmurD8qJ/DaxTclkP4+oQ6GUv7L8Jcx0oMMgX88z4c0u
1OjrFL6El/ze1HoSIAxTKKT2Kq+FXvy+hRn4FokYSodIPPkW6GI6MkBfxV5LoZpe
pz9YaVgjbSeZD8PfRCoJs/XQ4Y2c+T5dwmhXm1UBxEjqAo/I28oe050nkchzTY2b
H5xUv5/Ud7IKJTvyfHnPyLPAdUc+hP7B6wCd7debBzE5x31HB64FjnTH2KsENlmB
TP8Q+gr0Ey5CWLumj//upd5lDF+cHMbeDqetHbxFEYNa9ehOCItpkPX9hmksrOuN
wGA0ucWyZIM5Em62Is2TelR0KxDDu0SZr8kFQOHDq0k2/AfnpObhXh1yW5zwZdu1
rVhCORAwBaPmrGuuFocRUsJ/u9JbqdvHKJHgb4mlrR81h63Ia9ywzx0r4Wt/nKRl
/j6Ajxpwdtp7rdkYzION2VeNa9RCnZIXhriavQya+7YDXCTTpbqN5tkNWnM376OV
VxyNRDMSFGvg/Q3hov3rcbshHAUNqgXCHfRgZSHZMP1oo+v2enllj1xee8Gren+C
qvLkNH3SLEEJONT/uPuVip0be6F8OzJSXqcZ9JYDnjamqxR1o1YOZUz3O37TXr02
CBwmNPYVyvPtDBEerRmp73+Kpyr6MXZY+hyCLBwpbBuF2+/1I/kUDUdmVDCKX5sB
uS6Apt553RLAoz7XiSzH7J1V/+0OA8aw5TbeuTHAUJUTN3odN+xVkibtWSocSb65
8kmy43m2yK0MrXXkrBh8WF0KACS4d2+X41ZkfDoXyGiiZE0bP/CRNccz8BHQqhqH
7OfUrTcpqiZO74eG92aLlJfQ/UeD8trji3b9BADxNzxjIB8KTs4chdPYyckOpFyp
FImSrUuUpArdaq8q7YXJFwOiPUWndOzs+UIJnKyu+WFuQwn7Eycr5QO3ztN3OzjH
EfB5+V/wFbDBNdAs3XXHUzYO5L+voXCEpINpkNo4scrqx/i4OVffvUq73/3rzu2G
zIIenyl1XmxMDa1zipVNWLmDmoGjAP/2eLcodCJ3+cR4pBQwJYh/RgC7Ms2UHIGg
EBzBadgrR2KtKPcqRX1vM79NNTYCA1m/QKeAOGILzvfEYyGyUIzs1rdh4wJi4wEs
cwNCM4dGuzIbXJkot61GD1oZqowQdbOLkGig9D2bY+S+XFFWPLw+XvursBkodHcQ
nuUmuYnAwAcE/A/brTSDdoE8Vkm9CZ/iksbq6knB0xitKe+ys86bWBlLWd8N8vAY
UJgn+EkyRGbnazn0IrHZf9WTwAtatmv+7bs5fmxnJpT2F+zm5KwsT5ZreFEdk2Y4
QA3X+4VW8YwbBHL9ItgdJv2fSPqfd6aLTV7UigwvlkgFC/wjsVeaKy6CD1vYd3qf
rLUe/Jq1wnLEH1V8BKFgJJZexHlf+BsIC7LhsHj62WJgvROYuqLc2cNANbFSmq+m
zLPyWU3CC6Q580oaczOQoRvVGFQg+RH+Ua++mT2KUFo3F52GxUNOzZDRqtQ3b/+L
WFddt6XNknZMYOL2S+qAecGz4v9L1Q9ucVcvO4GnWz+kMGS5O60a3oY38il3MuMe
TKra8v/FFT8eCrnxthvD0EyPC7u/KexMkGzoDys13oBWg4N6j33Z5/QcsRSBEXuo
ILfk3eUCTF5h8D7iG2XwDhD0TRvVoy+Pa2MkWknBL+PSqD+0oIHQx8IqLbUloKNw
/xcCBFZO62B/JADyqhkc35FP3eo1A+nNX6zBfBc2cTc/t1S2vynpQTeoR0+7urQv
f4YgTLfKFPiCusFWiD8DUh5eWj7aLO91SrRsgmnfcyXD9A6yzh7+03qL2nCQJB+X
eX/fzlbmP6D0DtkDnlTzL5QLElJ+UJw95bsckNRUmw8Fi5/Pru6ecDiuwzCMT6yT
Ji5ZrXWlNvdrHsEzyOt3vA9/T2E1M616LerdvK6g64Wytozf8wA+6jM2B0SX+TBc
hId17mDS0kPAj0D8N3ysl0+k4YOHoBjug51z1AIpak30Uiuelt4Eg6kZUABe0Bbu
KBElcCQN24Js21ef0FlL6t7SLUHdk+Yz452uKSbQsWXXW8qXIH7zzlmkFalckx4r
8MVlNZjQLGxPHnSBICZqBIh6t4+leRMBgp3nhPbnFUYBUSrb1SwVtr31Ypq3nRCm
ot1XFUSTdWUalAusKoxv5V9zNeJ0ApqMXU3a5itirOrSUQ5SIycVj8Q6B3Levugu
VvNBm6JlxzX7HswbgnEHjy0ZKJ90djGmgGQJKgrNi9MUXtE4fle2gMmycVMm2xUH
DwhhZvu2/CzgmquVwnzxmZOqQtOrYPikiCIqETaxacT++vrNcPrXJyzn0TkMthz8
B7RvvOizJ4bPkYfAoA2EPwvGf974S7vkvPl9gvZY4ma2KITEdZJpsrLp77+/A5ZR
9W3PcYzxvmIKJSdtpvGQNBQrx6KmaRZ0kQNaUdy3SmoIqs1omNmOJtn+ulBk2M+D
T9UjW0VeB9trbbDCsZJCstirZuOSSaxEkVyS3ujLAhGaiiJtiZ31JmFWWlGS3GcB
9F5+Raq+cYcndCX4eAG2tUSRcTjjzugrWrgIe+e48oGLSgpgxmE7FJeuY72siIMN
6y260HFHEKgL80aHzPD77KU50XfODjysZ6zMBKgL8M2yRYWNqZR86mhH1RAwjh6n
GwCDupgP/0OQVz1Q0avBr3qxoZXsETy3vqojEqFgPeAFk6fpWHkBqSSFTNd28X+5
kOfWSO9FzJyBKQDGjXl+geKNo/imkw35pJajf8unJDhWcnrc93tx4KgpzIGf4SkX
AigB14/JsSAG6IxTeX/tQQw/JAFuZnx5QKwrrq8uGPPHiBUagiLOmcbC+8p5pvVt
TmLImiG6D6euosVk5L0PEZzIuzHtn1JYGpDBHPwvvE4SbGw2b0WG4IXvtQAz8D1U
cAZiDxEP7kA3OqYIYDnN1mW8906eiXk9C6AsAsaMF5gGJ5lvFlIHgx5G3SEQn7ZI
bjO1ho3rYLH3NmP7+abqhjsOlrOwoiNCN8iGW+Y1YLy2rSYWSAvIkJN13R3yDE5a
hec7876UqQI1mBicGGVQBAsA+HpPJgvTgD9xenLlyB4Bwh0DzMQz+/gJ1awciNO5
wDYndpacKN0KZz6Kg1GIXq1M/QpIS0aD7R2dscezC6gDR1FkHs61Z0tRMMlvu8Zm
eUAz3OvhcPQD0BtbvJi6R+KnmO3ItVpZ9hobZLbWBb6Ys3ajBbMWIh32RNhbUE0/
61VzfMXepXRpoLbs6ScRqwLN5o0cKbH+Mq3sbdCfOv8MJtJq6DjPzveuLehR7Hy3
JWCqw+wTcJuSKuCjMtrxjDsmJFw4dbCzkPWSEvE205Vnn5+i8GfIrGDLoef861qX
RdhX99Ipx/kcaa+pCQ36GxPnFhP82tB0mA0hi4bP3NDw9jm9t2ydLQlpKnJLy4Fb
6UCGkdVoiSPvejiIrlb9TgvJIA01W+oHwukQmkLgmz+P0Ou3vWiayQiM6E2QLVrN
k8tMem01SkbsbKH8Zy6rk2rkeUH31M2OrTgztbMDxiGOKV1RWv/kewUToNLdwvPR
w9/YizTWj4gTraplMCYQ7uVKw89AxorTWEdNoT/Kn7PyZf0PI5MNeYNNJhGQ38EB
8aGx1QqhZbiryKW9YhjPp2Q6Ix/DXCWkabjCb64FoA4YGRlEFRaLexOqCotNp0DP
KGl92I+acpE3Y9TG4A6VHnokM0lbua3ru0usW6jfLolMxvSdGLjPtKvE0pahUfm6
/PbGsybLsMncEfs0Q10tIMK7+REpQfZILWp5WZyRjs2w8gBpAX2jPWPncpi3CO3x
1IDw6NztvLp/WAYU+TeN0bgE97JJ8xY3DVMxxqxRIu7QY2F/gfiqRowZGe3nzoZx
6ksMUQWJFtvefwah15KxQ4mIIFuXLjUIdCMWgptczioBxaPbb058FbY93sU3vTUp
KI77xj/vzHwTIjCW4iDRnoN5Vq7YMKQ5AnZtPzLKcvHACxR7bnE7WNUKVZylXjkb
6O6ZrWHu8OlYRjKMVPRS+MiXJ3hSb7zFpynBTI1+LlTdk3zCSn1RRbdzCfHrJKxe
936k+PYRxbH0hPEJWm4cqhu/6EKoMbppmoxPfQ22IUd5dVSauUxB/75qAf/dlQx0
XB8d9jwBqPGa6I7sD7ekIa/MRV826He2rLVqxz7OTiNAPPxuKASHCqKcVhMn6guw
sQc9VCAzeB3bMZvqFMaLFTLwFUziBMDNPGvTN/WlbChDC+JhkztbAzjSas6QVK3K
puZWnhPoCW1TlLzdRdTgr323S//dg1Xgpwrp4HfecA6L8cCQbYUl2OvduYsIKapO
Q/K4FMJ6oDvb/OAHP7f5H5D4L38oAXD4C/3ITd+/j0zxMOiDgOFyDSoe7qODt9Db
/Oq7rUQbnM+OzrWr1H3Vkmfo2NpG3lqJtCt9RL2tTXOlOF41x3YF91L7u5fOrHLu
mcIkkB9SU7qfXgQD1jtyNwcrOdbz3MynOnPZTool9gjCEXaZ9hQdexfI+E1r9OHv
m0HV4ytuuegXt0yFbg8ImWI+vTZ13xNuo9uEQfK/mqyrPedWtWgoLrG4ZG8P9HCk
GfnNSZUnc1MGqPHMacWrFC6hPdYK3bGZ8AhY9NIqQUaMwobeI33X4MDRhwwlgVvg
SXhps2iLlX0/MqiG1qtKNoBd8ZYOkK6jeIZeYTHpxfV4eiyocvtl9CwgUzafWPs1
0yXxoF6bAkbB1YTsbA7wj0lv9tLgHbQGpSIZXDwjv6n3wgqvKp9EWnzxzr+IONWe
GpfLMaFHXztkkR7y2nxyEL+lYGTq1Ikez+/V1q1WwiTivuWHenTOid/EeaUzcz7E
aMVy0FRGibaM67WpsZk1onwRq3K1XQT/HB5H+oIppSHKnr6fnveg8K91wknGfCQj
Np9+oJOjJZmLa+KEBLpOLZGD5/cKqnn90HsxfJg9yn9ItCP7u63BwIIh2ERUSrM9
xTyxiaFUKLZNvmQjEf5nrcYdh7CZ7QwVIb+lYFL9przqWmld1rL+EzYCawRCAX5Z
z/zv7A5gRfZwSkiHqYzLIFffwjaw/6+0jVS53k60cjWOUviASdMRUFHeu0AjbZ1R
k7tx9qwXhdMvb4xRNi2ZWlzDPKjKs76k89R+dfs0mdvQlb3K3RwakEVKqyw1k5KQ
uEpr/1xeMbJwup87Z7Ua8S4gnf/+fPBRzYWSx8qCPR8QVTtmHGcWGYxxBAcvEj5A
LNOLmXTZ4X+rf0Q4u4EWcBNz0OIfJ0Z2g1J+wTsUPYRALnlVPeT3ZjYsv3eBqjIy
IVYAAqGY7pcNTNyycmfRD3kHB5NsEJO2UXEJ44mo7fYVumSJtxpQi7fnpfg8mx6C
kcZdm3lUc3NXYj8r8pzSIbhnzq/E912CO6h954RUuZmTDpQHGCa4REeFsTDqc/SU
i+QYMkFm571oCkaFpTrXQQtWkzg9AWLlwf8albspLPco+fpWNvl8BzHh1XvArIqh
eX+wHEFxkOFEaxKcfqxU6DZNOJc2ewLIKlV4REogKBXBgThpxJta8Mx6knqIyTTO
5UJzsGhcKrWkdZvL6XAiP1yPeAsj1SZ8QjJPqtnuCq66Elksm73lOPjVMFSFnMNE
TZvZtJqd9200pwxyMsxGREmY3t3jYTMZr60TL0N8M5Cehfm0FqfrvHtMwayr4a8L
EU+qcl+OiGwsdCY0uKSYxRGQ91yhrclYqFasaAFX7rcf7uUXpBheqd6yPvdKemfY
x2dmeMpulMoRdSW73tOkP2L2tz0dB1pUtIeUenG1htDXurpRbywVgtummwavxa7D
JJivcak7Mgf614WL6ZGtnZwKsmBc3A7QWKyl3YbWhqwvNyrtoqD/AlQG/4h+lkjX
rcEWdv0IIkgGHJaOP0W14T22HE6zgzgZ11Fcb/Q+TB16DtKIXS6/m2gEK77tCHKn
ERkJZoRcbdkwTsrmU3NE5CRgj5TLrn9y6hCbHjFg2GeCN82ACm+tN7xv9IyAhQ1C
Kg3qVoid8X5+y6zODUVngLj/SKFYjXAosTMq2OMtLYvorl6jffiKdM61HEnijI5o
oIFOvPCj2/GKjrwJmGqtUCTl83lkDUqkHjzH7b0FpyGvsMgJNCjvAFTnCE5ZUkuD
psuP0hg6DMzbbOnLcCq+LYrGCNbjdTDeJ/xx1A3VQmbWG5YmyHao7ZgEBkFb7eC5
BANZBP4CBV20t00jMNdMQ3BiuVOU4DNL7iyggEGGjTtIe11B5AdpdKQVg4JHpWml
4gsl33KcVvqEA3/hR6vQ2Ajs8z+QbEgBYkoq1hjNPrY6rMPKKlZ/ETdF6a/OcAz8
DNmzwJUYDOIRQVL7YDFPcC87An3naGUUDAsWV/99GZfleUydX0CfUeZN+0UZHAFY
XqbmemkgGzYtj8ImWd8BP+dsclGnbhrW5bcrWHYYI5Fm3k21i2TcQPzPNko8XwWb
L94xo3lMyry6KElIDBg5IDGT78bOczDZlwYttXLVliEU4YnUGceEeFs/MpCGIJ5z
HBGB2MoQ+e4vQVw3SJvYx+Mu6cGp+ZrHzbLA9G4uZ/MdUmXweXwNfC7yhBJDG2hC
+Sx3bN4v/CXLhowswBXUTLj7Gi/ukUsiefg+p9InrsmDH6lblWxEb8/60URTB+wL
SMWL0+oTGecoOOKBe3YUj9cJc1Wgjkw/VBzo1BK134lLzShhiwSBBmp+TyYf4FF4
3v13ArY1Gj+3n6auT0NmQSZxwiuBpIPXvfIjMmu0CZ7cHwlLdFbm//vQQyDiPHRj
5givTO/o6lu0ZGfncCO6Vk6Ff3Zf0T9SXxf+qKNXViNuYwP/p6lDoqDvZv17FAVV
BoudzL5q4GFEppv0pyf2qh9H1tZwLc1U5s269U25NXz7TQ+7wfQ3zLIFL6/Tz4fh
hRVvveSsPf01vL57ul+kKtK7IrHbLyl1Kw1nj06mhbHTOPGrVGpmhFY9Vj6PqrFf
wFng2g6qowCTr9e58f9AsCKpEFcmzWtgnXAsWK/a8YsRhESOXN/eGMOQYNchaaCy
W5ycy6kvbLK8omIPTooOxZ3k+sZbvtbQZKIECHvCGzel+w0FVe/lGCYAE7nEfBvx
AMT7PH5cYzpouEM5cMB01mBRxOrxQV6K3u7VnMiYbFsg+yQQvRlVnHwTPS2UV/AW
fy2QRB+1TmPbIaUO/9TnCvWfFLsK0IDIRZYXf7mvIzc158IKy2k2vazV4yyXBFUp
B4whvgHBx6XyzHjvU+KewY9bs42ETpVBRXO28lt2GAXAE+IOLk2zVF3KT9u1O8ib
IreFIhOMBp1QHlnDmjMx8sc6+ser9IzKpsJUdAVEfaxyNy0Hnn4J5tTHulxc7nly
fCsFBU5tu/TAQ1qmE1jCq7ga4ZOjfciA44P3mnBbhQ2bIZpX0Vw9WOfrMdG6lrSY
jeFkq7dTlcFIHHBwqXh2p5cuMSO28kLiQXn50DmfIqWFniG8QQbrLODe5OW7afMZ
sHfJ84BmFKaUrc2EjD5BJ/cSCn4UVmqow9nMCdo1rpSHZh9wOiL6qaVpe4+DcpmJ
OjI9uRHmoFzm/B5gbgWuHqA1gEMGZn9lz4NC1laVdwq1sYWtvzqQi5PRGq14LdOs
G/PYMGPljaR7KPXdtuK1mEfId+FWwjHntfbDAU+EPib/elVtC7LFqALvsTH2g3JX
wDxRe1GWUW8dibJjDB4O+u10txlyBH5JJ3tCf8xPqR3Je+jeVC/C97IZ4OspOjge
9buExqCOjGPI0SZ2Af0G5DGh8PftcXBXAmz176vVy2byzIbgA0/70VIDzmhkUbsx
Ds/u08VhS6XtkHkqLSGhTwNEF2di9fij8rySkpr2IVRriD1D2WqlrqyrhduEVJtV
BZa8+SNmrVufFQ9ca0pg5J0xfYr//VSErGsdfsBDlxvegcnVC6u58GT+tdMequ8y
Eq7WC5PVQ40o0ZLJJCBBNnnXOx6BjxWKYgr4QNCPS6Pth0/gA+mWC+hyXeucqILY
8+/02b6DFzW6sYkWvnO57jDbBnN20Ki1e6PN1biI5trbMut2FHMvXXnAm0+4RUUo
6G31JHMgaVIj9IYf3jjMa5lS25Iub/N95vXQpPQ/UeIXZjBhAF++7ZRv5WYD+Mpx
/PC/VYGBH+uIpNUg69c6sV6xRfT2paZ+Z2n18llVRLDWQfmlCN5/8YoXlhkelaaK
GIurMF4v4oXR6IXF9YeYEfTXmUtOCrvibplMtwdo65O7PuXhNIclhLL7izqyRjYS
ujFibWj9jXGrswx15BU/sUePk9m7Cit4aJof4BZgxQHle7Qq2HpMnoo4XN0b2Fzs
932dt404Sw/DgS0ClOXKhrwjJttkrich/1x0PqkQ4IoO9u4Jd6LmlLRc0wqsQWWg
6+TucAOfb73wNRguwz6ZYbcDouHcqjbXm3cRasVhj4bW71uAZpAWlyGQx6SO7zrO
rQ1Kq8ATSbwrG/vHZfl//B60yufMO1S1Ovh5GTUrPSbbQy9EYxfFObaA9/GWL7ur
l2DeAI+Sx5y3fZGzz7RPUnrH2B2UPOt2yX+biA3CsKniIAAYjd5I/KxJiovu0ujf
NXDZf4qEl7IYHn9c7yopqm+fOLl6BT8lV0g+u2RUQ/okyZvyz4sihboY1BfTJhoJ
4AoVv34Du1KqP+x0oHhVeYaXQedSe2GxrQ6HXSdoVaDKif5g4+NqkIaIhoDu9XUa
PmAtiN63+2u5C+PsEsglpBAEQ2d3zbWLTzYYP5a5EKMxeatyWKv7eGu0hNUQ4j+I
9HD5Fa5Hsp2+0h1qerHwKueiHPcRSAbU3lAY+ZPGxWrMYnMe+jUJRGXCBLOGn/sQ
HLa+PxZf+VpocneWwRV7AfVvUm8J3TCmh8bj9rGX4vTa6OfBXUP6JTlt3kWOPwlj
BopSlx/CtJuh8VDWmbH/mLIOZkewHrTMJFeD8CTMfbNRd9uU+7cQ1VHX98EDJiXY
ltbnb27Z6RPMi5/0lXWQoP+8jof9ItTpUZSWrI1sUmLITuzuVOQ5A21rOMrsmHQ0
CNTBssI7s5gQrA4SvGaZKJO9HysFoHvttAnm9ct3OkSZ/whTfErH6OGtSsszBYHC
rzZ+paujTKuQrPmOstFoIsRb3QioRue4NsqQklrw1GnbNAAJI4Jne+LTVk17rT40
0ZwQk+0rmb6IFxlV3SKsNdwKp2aZL3P1J2C22tpCPaW2RlZ6OxftHfEb51SOvhZ5
kLS4h9LoPKF5/CoTrIPNbn7QTlluCgSbL5zRWkPQydPRtCJlpiC+Ov2uhbZ5ye9X
PIHA46vMnNBcVw4NCMdXVpeo4ex4gY8VPfOzJdbQfs8pHw4KF4UAe7F08B8x+vAL
BMuyMiCzVqlFyK2x3uiOcD2RbMeVrh2BWmlkDVO8aQETV8cRM0UqOnUknvPElpts
0GM+Cjbh06AsnfBguu/6UINzDHu16t8BnXifOaF9yYgVcu8hfEctNBTkC6xhlmd1
BHdboTlS70CVsbTx/a6vfaoV0EVVrxzgD/r91RE//v4pbAVv90TxfofUme3lW5dl
dSSo1GBgcMCI84mqlz2oNLtUxxYdGMzgQd8NjXtWsH97hfpFpK+djSebZOQFmBiW
kVGRRIUBXK01QDSuC4/140QDcnw3S30hgt1zPBfI3BQfMhtlEOVx6VlU0XNyP35L
qvP9M8Sv8FH32NNFqoty9wyztYHXFCjNNNPq2mvLvWGpRiEdRr3UWoOyxiVCGAaj
C6TFG46QrZLxpuTsEplX1GK72YB940FNScPvijOgfp+NVq0I5ZsLZqWpNin2/vAa
UG6BJTQlLo1oEZPnseANBn+vYH+ixP3Sn98FocL+HofrPZn7aN23w2AVmbrizwMU
K92YdEILECTl8RjS0VxTm2hilHSme1t3HZEsM0WIYHyMLJWRXZLuxBJ8k8vReNov
s02Vr+ouqkatabWcl6bPUJME6YPVxSEEc2Rc4eKki0axWF4n5dI3ujuHPI8neQZO
+xbpUOuHNDG504uvnxNJvQjZtfpJ3P4Qm5coSSp3jJC/uP+FpjlarxkldswXhZgA
mc37cpOxCThi2TD2d/DZmU+onLVSZ07uSXOFwqr3mIfPpagq8gH/Bym6l1pBLgjz
UB74MfNvw4ArP5qv4JRlqK/aZa3smy/2v2kBVEFfIpag4dKoZsRsxgH6Ojvfnrvh
nl+YsbODFhv+xwGiyXkSuh92fBIhZmkJ9o6Kd7RiPtoZZ7A4mrMtl1hZ99Zd+0xq
WPkqdym3u3RPmw7qy9pxEXI2arm3yGTVOBY+YEG4hlIdsYc5zGz5ZGx7bUeynu8q
txPotanDnN9SNQz+RatAg8rYBsni3xxWmem9+wPDjt3WG/BA+POX6KXD2RUDB/ES
14Qqzo6krjTvCPHU2e9jS/tQIv+SLha+fbpm4PyMSKjgyQGIsD/SzJ/PAKa0Bd4c
XZqKz1L4qM15HovpSdaBaLGAiUzBB6uQIjs0X7Yj7y1a0/JAlvQIiJORYATM7NYW
Jrr3JjVKKU/hveEgZfXnv8tz1R+lbJQpcZNLhavIn1P/LuAn/1ByTiTjzY/POL2h
Ga6FlC+zONalZYglQY4OzBNFsFMIlS2vGDpSSuBggbuvEkYkt+qIu84/Yi1rhSA+
Po5tgCOkPMC3qS6w78OHkBnYuUr1fULtgL5r/h7M1NOEOpTvZ34VG3Hohvx3mLN6
hr/A7LEawsFSwhF3VykfVfZxadB0s4uJwyfkFTx/IJEwWb+5nLnrBKkoNn9QSQ6N
thHP3dGw00qeYP+vrQJUzHmZYydf+kB3z/6PFJIJxK//Qcml95HRHxuVxTF50usv
xdGknIynXCcCS9w9bQ29lXvDe32S2ZZG34RKwaum8c06bCCcDn1kWpDhZts9vfeE
YKn3HNVtwFydBR1tFAccwJCBzeU6YZMSFBISGaIJR4MVz/5WnUUWduB7qBzjE2sb
wS2CGuVuOqwnfdf/uTFXtUju1egmV3InGB2cO4HykcNqKdJtNzxw9OCmAq+T3Eez
ZD8PMNAzxbm9PXju7F+YSEQH+bHAhC76ST5t4fzkxvFro2viwy47U+Lz6IhFVfLv
8d3D2c87ySONGx6fV08R9vW15CfpBci292tf3oeBMl+RSuxUoSA/tNi6cpbDD6AP
Qe+V5k5/3+MseRYQzuRD1O3b0L5+brUOiMO93g30kZMCHruJeafTHVt+IuTJAzCy
JumGa/zAC6FaiqwEkO1T0DZCzecluJlNf/fsyuLFV34yulP6O8r8LdmvYqZEhIvX
2raLeT1PDBWcsh1eoLjf4u53URRu2nZsjdSZDbBA9eLo34E7IGvwOw6yv0KYauoi
NanpQx6FBjt2NywvQRIEtiHVfQqpmuv3qAOgxmw6UV5pwpLUbuAFZX0zyHofUi4j
xTV86pKUv5geoSM8NW3YVfcD+FmCvVcEThF+CllgW5eP5CNGYxdoEJkGTs2ChhHf
+dud2PQe/2ObOfw2w1VxYEBRkGlRuF/HR3ONmT2zuAMrVMg9nqxAXZ4XPDkdhaik
rjafd4zV/4a4D1LrxcVWiLZoEeCKvth16qSj/+aWfMqKgFH8ShSm2RzOEwpKBMz1
bt/6BppdTC25BHyvAC7tO/mMg4dgvTdCBEC7oCE+QM1FYxQ3MZKvMJQDyG/4IhCA
FUVR+aEsCTACFx1jhXI4Wgho73Ffd6AmaPYPbKSaPida8/0EtsNtZ4CVb584NMtD
m3Zl1DC8NcWvCahpn9umq9mNxAUi+ouvAK7wN5os+l2d1RwEVYF0si2qYbmAYZwo
IkjzaizZGsoRd6nMzLIFu6xZhcZgW/9cyvTtOxBqSV8v89L5g5UZwThcQcslBXaU
oTEQIxYOGHPI99sZz35UOWow7bAiNHBr1Q1RK89VpqNBVbAa6z/wPw8g9c+ZvDgp
rYO5uw5YPyfXjp+jfdnMssLpYotVX33vEBD5RO473Rj4CYiUnsl8PD3jyAERScGs
ljMaVh4Edb4hXiNgj44hIgopVBDVKse4GArVXOCW6COMplayMG3YTweT8ACP8CwL
HpApjKlreY7zyrUBb+vBZX16DHgRon4cGHJHUBUViOGQry0wBluKpm2MTMk3LMuq
AryPZJKYZqZ8yRINHmr1S+nFLXjLmfCo2kJWwWhZ9N2EieRRAUYQg5rI2Z/CCsrC
4kscVL1A5G6PuW0afkIV+jGJ24oOm98L0HHDHatEbiv0+VBwryGa2ZfFPkXbEnMH
cUrFE2hYwUgFadu6JtTXjJP8167SBmb1uzAtZsuNUvtNTu5snvq5clA7yXwDQg8t
j12PKX2R2MDfNyQkPmRrO5YeW/gRKMc6Km+/01lYcv/ZGufFN6iDcL3k9WZIqtGA
VH6MeVBhKU3le5gPVcVr3y+RLZulj9zSMf9cygPLrCVQMDURCm1iw2e6SSoswO+/
/Qe1C8mweSdLcCm4M5pUhRFuXiYsC0knC1PLlhxZxLOkCM45diER/OTxUJtsFraS
elPEBCiiB6muBtNHjHxWKzchWHCzIbU5b5wmbwjUR21ZkA79FYzG2Rhon2z08pFE
xbvFb7Nm/67kVMebCQFxpEpNXsMuZgghiWQJ5Zcgtb00jZqwnZiw46ilULolRs9s
Wt6C6CMZyKmaTHNyW2ggDwbslJj03yh0uFcxtZ0mXnaTNI1f4hTC1Cl9XzlNzN55
e3eq9xDr5UIXYX0jVz4Idc8Jxo7GTZ7xLO0qBmkHTBhb+mjPDGRatQQZ646jvyYD
YfShuHXfFYJbJef6dQrOhEbmd6halGSVGo2CsWis4IWoZeNCy3hRaghBdOh9Ti4j
UdEvanMGVLLc/jrt07TXz1l1eySJaXtoPQY4krFFUSdvJinYL19kZ1MPUfCDMVSU
B8BItbZdkVedUD5/OqrCl1+hgYVikSkIFMFGzWUhHZOaPFMuVbUXx5tkKzi5EQgb
bzmb/TyuzAYRlaIP9WRTLoIo9M5yWnU2HQEND16AXBxwuJ1gXuIP3UPBIxCvScin
kKvjTZ45ZvbArkpRMqEDZFS/wiG941dEEZ1qDv9fUqyBaQ0Zu5nT7CsZQoMRS03P
7h/67rtjr63PyIVToqM4LNKwGmuCL/tLjYyQH724MfnCOmVTJHhV7VDtSjQPhhiY
j+rh3SHCI2YwrifM5Am32QLiZUWRgS9Hlhb3Vc8+Fs+AHLxAbuH5/8d6Q4AcgCNL
kkhk2SNmZpn35oxUbaevYXK3JTnKTJ86wpf3Laj40H7efpeCchQlS/J9pQpu7lOA
Akr/flCufZHleiYCyOBogl+gbz+sQAzrsfBHwJ/QMItl5kdxY03timmmEvZWHIYj
cXNgAFiM3b9ZYduXx2jNwHyIwR0yMU3X3nKG/i2deazFag6N4FCUHsK9LOJYz/D9
uXXAG0HcchUJWpXN3wG47Dq87JoWifFejm3doWe5yGprjOCcitsDOz6zt85oGSi5
2E6uuagkdEEDvQEHyFD+ve6TGbA7QsDSnCQ7UEQcrPNlU/2UnCsHHY3KXZvTF3c+
RAdtJ0Ors5NaxR12aoOy7fP4gWTf43z90zHnwEUUKatKFw8JXSWAd6GDbQpB7GZQ
VbbRCSRL2zjQNqLFiQ1x9lgoIf2I99+SJmdBvz92vKCLBZPKeUcBHxXNrMPTAleU
lATMH1V87WfsN/CcaqagkdmD2tASfo5y+yak7xK7IrgbsuesIYmXVCkh+0xdB4s7
GV80V18p8uJfpkOFXwiqSubU1614JwMIJZkSYYhbfXRDFtvNpaYxFlzFD0U/b5AJ
DoJPoXcGkJmaDqLA3L012uBu37ai2oEDHbMWPi0l0ygdBxIaxFhFWwzWmXTLqBNF
Sfz+xiW1xsfQFk2p/VLTTJyR2Q12M7PYwRoPrD3xz3xvUAI+vqX/mIUT16+1CE3C
yKusmQWRwO6aOMdDTrvt7BzMYI6C6aC2fYIhy2A8rggi7maZHCRFpBsTRyHw9ved
pCa6CUnRWDkh+qVFLkY8jw7U4y3Hv8meQW8kJQEoHFbMTQRvy1XE/9XUPbKT5B8G
/aUd2bkvrWASnlOipI4DLvuhiOm+TRY4z8vwyOQQ/85Jizj2UdDx1HVhsCT/ZiEI
9MCSI5mxztauiZe8sMFNfZI1tkFeLH2PZUwPjW+qusa5faTgioJuoY+y40lqQk97
S8RV+DWJlBPwU0bloeaW3gsST75F+3hZhf5IQCFBySlDwobp8/YpWmbqIQPSQhwQ
Rrp8cNwS7GA228jgaeQlh/qDnEy644Ko7m2MJMCHIz9+vl7LbgZP7rHpygUBX1uN
EFgGpaqwjy7oHwKKE0stTaDafohW0KzUq7dqx6dG7lrv+SVFYmVFKKhg8cS/Ptkz
uLYVVTJTSKZMl4JGmH0hVKXloWsP5a7pt68vuCEZKJmJf2we7LnZZ4Da+JLDeQlN
sx9b7Nc+FhRu3jT/+cvopayvqXnzbUBSwMMhgs+0bXwHEOyXw6xhHHVCNzMo69bC
vepdBZrl/MF4qli674BgfVnt+OUPs+VayuR1uOwI4ySZKO/GTKbIa0dI0+f6jfsI
anJqU8LCwmb3pdPbC1VqGSiaaracbyRqEtGr+VEJSO/477fM73O8tOxERQ0Trde6
Mx0VFL85Q0gybrm+Bb2D5RRR2JHMzvUop2Yu3MOq07BLzBaydQbrwNus8j3qaYg0
IXdACMlM0xz1dbf5b8MBwY39gdtI3U1tu7L9QA3UnGHghoO0yzb8hKoaKNWb6d32
vSUKLMC+8wsHOVJVfpfs391YkhReqcoUOLBtWhGkeZ9ACxUAYiVufvM6LfXTUs1V
YkytkbndLhFtwIFMsGFfkqQrnEVxRbrowfGr6rmKXpnfTAG/0jUYscxZjbfNfJVX
pDG9jag+lNl6A5boMTputRJSxra3+ixXbTKhgTS7cAq7xU3NjT6WvqBAnPfxLQbI
+LX8LFV9K+5gGXiaez11HR3sR5I4bEVhTGcSnhv0onzf1gZic8nuaE06SwIpBuFw
feYyN6/4LeM9Yqh2BDMuX/zMwf00wR3pxsArxf0cgV5WBC+jkKW0oKZ7epKuUsN/
VqI2/Zi71AmKSXcYzC4FVjbtuTHKe1qYduD/nUoqh/o7iJrJYc0f8PSV9bsD62zJ
HQgfiR5GlSR0YjQf5p9J9x648yPvWaf3X4FijVge0ndKirYn5CFdxeyWLbqG5/+6
zN8vwwhlmOXWyu+ZNbuenaxW3qyyGhmgO9pudIJhZp074Hvs9448U9m0dyhFkkpu
6IUMX+YcmUufIKRVDjXmnD5GCO/jDWWbNcJSeUZUXliURxRVmNzgr6Pk75hT9Mmt
eCyJxQ3mlWA1h3ZEzxCdUEPMOgYRGqnXIzA8OpQ8Em7KvHJFrwJ9rug9X6a5l/+a
IRkO0zEaccmpok7kjzQWxQ0btCFKf6H3ivmB09DLKInxSmIQjAjAQjh8i5qOnaBS
tn9SC/c33sUvpzgUBWiR01Jn30EUtoYxT7X6A3Iah7zXacyuOyzkTZESi3OAp8St
4spd6wkBN+f1Wes7YwPnO27YKUN1rfdoVQmWR/9gLupaAy0yCquc2A2k/92O+diV
6xzRnXqTIudX+2K4EiNvrXJhOMk+wLzZ9iMN+H0Qq/rbKK2W24VEspDHzzFqqVII
2PQDivrxB8XtAnr3YVQz6tI0BoHjPYBD+rHB2Sb0jFTRynci/BD5nZq4JRMhzK/b
HSHOZMsQ8y1KjPDOKcy7lW9jLCEbq9seIKDA+AMXzBufJMgLY2TuXAiDf914TtBl
un74o1WWCSkB9rXFaNadGhtagoDEAWL5P4J2uTY7jKMxMFYii79n/Cq2l14qNZCK
EuRXADIS8WuCbC8333lqFlbasczRqC6FoWvyKFt+tjHWk6fnGujLGtH2OST1TY1o
Qz+DXwqQTwPHGlV2NxQI8BDHefD5pb0BGPOfTT2WP6cIoh0/eP2n5HlVISgs6cLL
XYOToJYlvrWbWwOUHOX1AXhAdmvqxn2pgsUAsYR7mdZi8aynKaZOyuXCxkwruWsN
EJyzMiRilk41KXaZmC7YYIcz7P1V9W/voaQCtripbm6Difu/fL9/NAk4tSWRv+51
zsdShdNSjPOr18Ajp/i/orEtSs1W+F5u5iJdW5q4suBT0Z+KoE57MDxUthqqIBWU
CJBz9eujBcdiITj4F7vteW1x85flqKu4fn1QnnRHy3pM1xrc3QCw1SK8czqVzfnP
YCs2E/V6BI2m6k3IRoOap0z+yrBigS5w3PQhnZU1vjJH+wnGgkatcezgbz/GMY/m
ogKmHaAIsDR533zb9HD3Ig0easVpKqoI/DURbwzSQv4hdiejWyBB/Yui1wLW8m03
Oe7j0QCtldO8Tn6TxUzPYEtq3wmXubYihg1wqQHi71c0vbmm7de6+OTdOEABbmB8
WEm5cZwb7WjcplPMMo0ALCyGf67ga7NBW0AoKb+6LyQWA+6uGFY3ZvD0VXI0AWLk
7sgHhMVNiWmgQfy94vh3ZCKz64rTtrnmekPxQbDeykqU0kBi7s91PNvD3tIxRp3f
8P0SJCevW8/ij32l1O87ZDTBJB18USLtPvEr/wWzqq3u4ZeCSSYkZMEVKoQw7H4B
O5HUxwgkccSrRMOPtDEHxPv+2kWNd0ncTD/EdSUWVBp+zyNPefitFX80InskkgzS
IuBd754+DFpGdemDwFafChtGV59BVCiM2OpKMKpTVq/vg53d7Jb0H5sJdEKeFvu2
bFH8SyKdb60cOs51+ZGTVzUp4o371iFKm6ZbASoFsd/1NQN0CqgyuzzuMJyKtqIx
G2OE9QJOcbMbVy9NPEP5U/Psx3QAgHjZaf4VfrGHAbkZ10DBIgi+xQgYUmozXWiw
i57O6rvvL0FretDvCIfQuDbT+DXXcpi9DElH7+9yEj/KcHh1wCJUaRvhC0SLBb12
CKz9vRpYVZQgRH/K7f2FcdrNWBugE8GofncmQw9HGeCE3/C8yX1Q2xpFrdx1yyVm
hTWD2O3riOTJ0aWz2tduep2lvjd41GKsubYYl0xB7nFP/Q7hcnBjRvv2jpi2Ot/f
xOQYlShAu4RWBSylaJCyWCxxEB3Xjcghen4+y8bgoFSYaUIwJS1RJwJidCASsMjX
6vnI97H4Gpw4caRwR6LG5umH3IuCvoD1D/AYhOY06q0QngQYTG93pj8YemPTQu6f
LgZwCXLWvYkXKh6pUAS5EezEG5uDSM1/p4+RxFvOT60RelsN2X5cO4jyz4O/HQgS
BDG2FZBUtGzJA+cwHlD/+EexFeVHnbqPiawW434dED+E9LUdmu/344VAY8ON/hCW
L2zWCmLoBgGcbqdiTsz7uucpqFn6jhXs2ZY41+GVJO5SJy39wPEJak6sjL9W3Tuv
iTJTRdvQdZUEOBz3t+T0hCNX1yOQufR4KLb6zE5ADlSg5o02rRKTH/YOuJzXDk+p
EMUn9M2y8hknWPufhGiZ4KzcoOJAlGv8o54pNQq3gE3j52IEsJjqrkNv/6Avc7mA
Nj6YP5CmcMSUVVnciMi6l2MgIGAkSOrR+2PHkiMIBguYkAvK/4r5stMH+x3MdHqJ
wLGnFpp8Nl3BLpYuwh/m4WRiWkdmSq2ZvEXY/0+481VKVh1woAcVYzHflJRB+HOe
JLlnzceyfUnHahPA3f4AhkuibcQr+eLuVc/RlrRpJxeLA+cWj07b6ngrLHGDRpJ+
1Ha4ClctYbbf1ZjZQpbja5A/9hsRKcqQ+gvIWJpS8qeKPK99XP26M1MvmAbF35up
PXzKnLuHoOnVhnihTJnnIlyRRKE8YMj0dKeOBMeOo4S87FAAlbmMjrhfNg19xtPC
jSlLSzdJ7wZ1T9pCDIN/mgvsezmMkUSyZimG6w6UO+/LeggHYOqGE5/YFRU5eWDc
TM6GrIaotS4HpceeiJUn39ihXfFnCWYvuaE/1Tm4Gsp6IHSqtAFgGjfWpnAOW9j5
cgmH6eiMW7dgDQV+luTtwJPfdLL9dRMPYF3E0/MgRWPVnVYr1BfybbeId72zSMsk
10y2KcDWAV5bmhUFjUiJ4ro5PLJYQZ2UgXdwAFb+jQHBFwD8weeusKvkApgiFeQJ
I8kDKAuidt3faUSBj/f9jmIeaSckWAO7s5zVijTo6Mt+47AjcKi1izZbwKRO1yoi
G8PdapiVhBHKzwjYc/+nzHj4JzM5fNNUDJPcN0TaUuCnYb7aIepLJ5KBnXBkEJHv
8VsTTjiiI54h//4PD3AFBq7KAYYamQehFz5UI1YSbBQZBnnBUuqnk+kUi4Gu7kmR
JJuUW9uOXLqJf6ZTz/iyMH2ujzsscOxCcwVapl/ufMjaMFv90JohiWSMeebmzyDS
cVOHKvVMDy6gLSgO4lHircM8eQvw3haxrDn+a142+/3Z/ptfp9d97o+GuPbJG47P
4hFio/v8FR5bAE/bpAGxhaGeEk+I2hT6KtZI20Z9+P9eYsUY0YJV8c2Z2/OMnQu4
pa3haBY+ue/NB/dxz2pcjO76kooLZRWfnN/lPleuby3n06EqIpjo3cikDeJ/TMDB
isBOJy7D+KRyYaMU3uN7yT1j3qIBjKiWpF+SjKqQldYkSFcv1NI3F2MOV8TZesMS
HmXp7Rm1sAgUNMxL4rjD3hKqf95Q09f5qPG6Iscvg7bOFI1AEVVh4VwxQmP0R53t
lI5Wp58SGLIVxs4YQzOWqwccequiV5ISNBVDJFj9vXgGSx2TV/inxux4lFsp1yp1
Dus3TjLVaH9czzZucrovZNqs4Mp8dFEpsz5/ak+APTRN9vQ4YcToI3FsYqv9X/3E
+1gScRxDnKdifVDFyha/dcr00H04WQELe8FaowP0gMyRArcMZ2rZt65nW2y5y2Sc
mwLlZN3Riet7Hz/A6K6WpwMekfhZawEbaaYzL4vGlrXnR3hd7M6meogKoQWAVBm8
oWLNYThG3tnYtxCTmo2RlcP6A35oVc+KwLSnPZwtxunvB/jXLPRDzUUs2JZseO+h
VZle7ZcSSpYQaC4TAbA/mYQQDCrRvhDJpetjQAEVNTVc+M7in3Ha6e6b7/Vz+dYr
ClRr3YgsaHjM8uyHvJa0qa/esQqznEW+wFmRAUNRiABzPEqit4AydNjRyp/Mui9T
ha64eFgSzScUmMbhGtMnC3qbGW9k0zMT6GqOX324h9Djeo86r1iCzhvgmyCgD6bv
Ofb5S5WVJRtbClrrn7jH2PZCXEVCH5RoE7vIn+ZbZSuXaKaTHseHz7KizfFHYIcr
8FohrKYn9NGkQDe+If+6mA/EbHZX1WZj3UfYLeGBdBgHtsqbFXkn7eH3rsuzY1Ik
XSMUfh4k+Yjf+GJneTkgGceiGPrAWAdUxTl/z5N1S/rNJnmbuFF8bFoCEhDDfXOQ
k6f2Q/ZzKh8+pAJ7EowWAqfX2ah7sJltSnjw901IJiRpGaZFt9unOXXcwa+FzSJ1
nKm5rzKGmTF8tWtDPRChSnqYJUpiTkjNNieZ53ZxFmvOcZRwMDvjYliJ9huLRjdG
DGFA+2Hdfd6E3X84qpiwQ6O+ifJj53fCXkbTBQUvdDDLNlXpSy1qDFXuk5xVM4e5
0cDhaLJdCPxZTdNnbzw75TKniQqJJYHmcBBCxekORJJoLsSyyUavqMTCMWrxwAtY
ThnudtQQn7lgmIMrPZx1y5cLenIJbYW7suGIFMoN2gIvctDeJrYAnXcDoGx4tSAN
zaknJkxMs16Cj0HMbrCby7jMZbNNOuClo5S2oVoHhovC6tX8WC2kbam0hf3syljB
CyKZWYu2LAWQsy8dGCjiYtASaTmTXvK/Pq7YuENaLH8zasuLgzpKQaZJ/8lI8PK9
ofHKYHYWaXQiJEqFkYPwqVZjVcKb3r92tPlsNKwaT9W78Anyq4u/kCiy6VmWM9d3
yQOeNKMeHFTOlp6Ce9myvrfUH/APb5th8xAwqbcuZ6hUGaQYaaakMtgZySMNLgM3
CKpgrPxBFZ8FTnqG1qmnXgBYrf+IbAVy6fboOLcneG5uj6/w+Xyyck7di5BO5SWg
hukB3ENofXacn/sxZNxJrzeyu1XRs9nw9Pa1OAvvB9WKie/+9z9wXXw69yfC/xmh
l+jZDIAWgR8mY0n/Yrwu7+KFL09fqPPekISh+exc0wrV48nzsqiyHYY1q8E+guCg
MAsbhK/3ZlvfvRa2QUhVEWPr96pBjUheqAziqB9FJNTOonfGugCVlkXs+H5Ckjc0
Yu54Y+XCwvR5/wtTH9eTa/2agLhXqWN1mzHgQjhPMtlqWDM2O4fFE69Uoyhshp24
0MJeqI6ecaxovs3kVNRO7pGMQOOLLuSSPItM3aGzFEtgcKpLUcSg1IHZ9RQoZA5r
uHyEpCzhrNo1YRcA1+zhBqyj9mnZ0Ste3LM5BXTsLsYr+iHxoehxpueebMxnzNxF
WzeuEpWblnpRvjRg3NCNAbVhNSJ3q4cramuv2ZD/m/fDDxQwlEfSpESURiVo0ccI
/VJHIzPcMHlj8iaPg2QTgSXAmLY/+LWjP4M98QnOeuyup9fuTHt57vSiNzKekHNz
kb8W4f04ehX/38gMoU/o2XBIFuAA3Ip5Ghznc8hsFHqBgesyly2nmF+UUgMpQBxu
ZHKCw409ZoDllBZrdTlSGclkQRIccPipHRj6oN/0dRaxf0dOPE+oWj4Z5mmSMwwG
77cD+aQm2XsvJ6lDCGuBwS9mi2ztVSpTNQS9zD8CIf1my0gjvkPxUh435SXMcZkZ
6ubthSzCIuJ+5RY4SZ2NuuP4r4jU7kd8Ez4qQUFGczA75RG59OaaedUhkk2vgS+P
muYCdk7SBBAkg/Mw+9lGdKtiV3GER6Bifa2G/y9/hvG58GAUr+ogTZCslTbxCwOn
UHX8PoO+GZwr9rpqCtta/JohFr+t/+26Bd8i6dvPUmFtbgsv/+aEikR0xKBPBd79
Pnu+5io2jf7j2sYoImAR2pOXQY6lLoZNkQNmm1lwB4FgfmH9PQORwr+kw3h/Uklz
AInQDjw4Fy2Odhci9oD90z0KyS7rfwdy+OVfVnpxfdy94J5a3N5EQNRjN9qH3sXA
peHmBSHqpFbn83vuuw6GyayEHXoycZTo8o43EsGyhqLAOvY4gPXy8pSpQyLWDXBJ
Gu9m77TpWcvT0cH6jwkfYXjGcMUGxZ+zslS/0hlLEK5TtFH3UH8ben6Xa/GaamXn
7p17KRcMdJtViHtB1FlUWTAk5iKihf9D8p6NtzqZBipL/3jYUC81H6bZLRDCIPm0
In6d0oBNdaAcE2yAU8kOsWVlqH7uHLoJym+vWCNbqYwoKLUR2J+H+bNB8KbDdMP9
Ez35djgGMo+WEjSxDzwjO6ltig/ZP7DkPEm5DQhYIo55oY22KJUkU7kRY4SrmqU4
MsqVK6Z4RjXfkepCr858U4qnE57g6llIahQanwE3zHb+sq2FBHlMPvUHKzmaKZtK
FWwaPDsLVAGHgR5xmnVZzMNH169xLjcuKnti4erbm5KzYTWKtLR+gZsdM9tPloz3
n14FeSbSt4BWwvJYA1hmEibkUDhd4FxCvjWQ/IGiZsYa3OWKMULe8XK/k+THFNSf
uQlYcUd9jsbRfFevY+sOlikm+OnuTLn2zs55imKlpkJD5GE+h8hLi1k4030iFnEP
ivh1gghCHsgjrEFojP6uFD3CjCUkPyQ1vp1EbLK+QKTa77D3bSYXPxS13gmR2hy1
Tvj+9/iDvCe2iPIjM76tz0IQmssjiwKxKj0CJqGr6GL0z4zo1K1kVVC0UNwgVBrq
JvC6zin1wQ9ixQm6flkHGMmkYNnewsPYEQxHzbeq6D9g/a4fxnPqbHwm3GaSh9Gz
UF0wyIC7K4DEUicUX4bTUTPCdZqQPjGrpaBXehbcaWke6SmTNPFzONQh8w8tTx34
epK1+WA+zxs7oWBrSRBpBWUYo5RruvRWNpCihqV3TU1gWLrXmqvSpbq+HRpOBmiF
96beB27ENNUFmULx294IsmqqxQNJf0AcPigxa1D5XDc5baYDoCXv5LS/GqYJlfE8
F7R7sy/KhDWmVEFfU71H1vL1kklFCiGsU+kW1dBo94js9ycr2jl9TZ46YfnH/qPg
FBHNYHasPvnaoKipWS4eWDTBThyvKN6N2qe42HpWtWQjK5vQUUMN+KiNDqNhmT68
kQ5efPyewsDSeGPdwFocdxJTZeFv2gAzcJbxC3379tsL3oAfaQ0OgCxqyTX0S7Oe
bqBviuJNPDlahk+x0EM2dypZpTp1xDQYMejRsyl8l4nwG5RT414ceQxePQ2ak90D
ElxO+5m1xACj6QPbBecAGqah/sB2UDHRGSgcRrr+U5uJWq+TMHBvLrs4LP7UosQI
SK0Oko+VHHl2YOJvOQXjJkJpyW3W51nxnLwGbskiXT8OnDnjNBVwbaRhSGlUE1ch
K4ISkYKfB7GXiEVatpzcgGUIEw9BdO2xb+HwIOWFq4TYldO5WJfra8P8ySO6fRrZ
5J+cagsNAjNQCYAHBeeco5PzaneuE2pwvP5sNCAR09IBVIi1ApDFwaOUvZUzSGLC
eu8fwCtISCgI5wwCmkO+gQIRwX3fUffxPLeh0L1SOKxge378Ay+ijb4ggLxyDFdr
S4rbR/Lu3dyMgGXh8JlJU/0a1EPceZeSskgu0EUWbiD6HvIzBD9Gj0g/1bohBLWm
HpzGM6D9UNDp/K6nBVjlemdhBtCfb1+pRE2JmCwu1I1UfvZExYqHDmueFW3DOkXy
zmM9w2EWIFLOR8L4rj+Uj3z/UdiYLH/SNMgWtXCh3qTuwrTqSuIBvPcputQ2Wu4f
Z8U7FBz/w1okLaAu+amyl91f3xakbFACv1oH7wbhLEml2GsFMdY6IdvOB9aYRqYS
HCpvhe++c0jRHQWnOzjVq3iiAWi9fwD9iGmvxkO9fa+bHQBhm+0BcdhUxfSbPyCG
HJkMUxYV90JEbuqUr/bkavEKia58MmaqttMrEc34PhdHQhR5w8fH7hnrmDsId8Nn
PDuah9963sF5LjQnWJVU1IgEx4ol07eJg6bwg4jMYlZQeyyxxrpIAcdbNDXZjKOt
kgSckdLwQITlhU2wRMTLv9bhda2oo5A1mVdG+YmGRi9S5yAKp4SvRgEutLoYTRQr
H1kxXoCIhDhQgSCaFVHD1nBNH1IgefisWKYSDrjfctw8PJiWnpVRPiVLfm53xO8q
KUSkoCj8GWc6geqYjj38KEFIpymEnMyXPIoAi4xW3I0c11mOkhtiD8qyHp2hBwlU
FXWk8qD187ZzkMvYhyFHoP9Y4dZfCBA2CNRGlqKmzv5xBIomwkdweFL0S6q8YWeJ
m8VP3BSpF0Q478tWL0TP4OAaQLOxR6WvYiFP058Pnykz1NRZPtMcuoJ8jHbIBrEc
SRRu+xrnF4MoZGKAL1IserN2PnZt3Z76OcbiitGXN6S8S9xtdbOLklFHswX8PaKy
krz1gYN3+OeWCxdQMKS81q/xc42TDtSv5sAhMlKJzXQk3VCcWHuNbZ+MmpuKOUNw
7R1w+O5vzB7GeNycm2u0N8kjBJ8evJy0biV5hcEg0Yhue6zJMDi0tPA+iJwbu3KK
bP58N3q7VHPCL1Rr0ae7cdx1wHTx4lmlS0A4DFfjnQNIrylFhfQTJlgO8nD8kKtB
jUaQ1xl+tCL3U2Wm4fuaPhE9/+RBUCNMsKkOaikU348+GDO1x3lgfarCpxO+I+ph
QbMpNBadYuf6SMKpD9cibv4IaR3ql2T1gY9WPss8/UhdRB6ddQcQyz4h66j5FiHr
mX9f6o4U7hPzwZPW4nHEnHOcgT3TUDvqVTfFzsZHvVIOr9GgQWKK6wsfWM12IOMX
XjfJ9XmohHzOUS5X8MOIN0VWNmBZs9vkuxH9mreYLHPPjgbiY/4xm0/1QJAn1oa+
sys9v0if48uWnFnqc22AKZS3RitFuXGsJCLw726kP8jIBKF9np6AawSFitN2L3Dy
I1Uo8rdivciRw8SBMeCfAp3ankcVK2FQ2g4I92sh/TYc//sht2PheJIjRl5OlcPJ
+N+V+UYNrn7PprZt9iCCHfVKH8DyuSt/CVCMtQOspZWMAb/iPuRMCgiHEYaN6YbG
Zj6B6r/cEaqPmNmxKiEgtIi9zlUJ3ZpbeiU1p5ohsDmuRZU+AJjaIHYMKuu1QmlT
vzLhuGR56m0nuIZluWPQDf4DreJWrExCWbry1rMM84o7xLo16aLy7weq3loYLfBK
sW2SNXDbR/9bhCwDq4T+4X+YFCJGmej9zSTXD34Wb0XG6QPKv5YRmGiATQ5vX6Q9
yk7hB+YUpJbPItFJW2yI+0Fc9fuXSTP9wJPpRrhuLWCB6+VQ/DYZmkSx5wlyWtaM
DWnhvancbBWTEVHzMZ9fNCknlaqs7HlRZLSMXuP9hvhuXH/Ad4rzz2lnHYGTz8nh
LdsYV07fjQ8Jm0piIyD3fjpYzY9FoDlb3Dsaj7AKMxW46as/I3wNmlcGEin6U7sP
w/PfnjA4hmaKBtSFqLTPNpcrqAZ+m/iNzkSyH0gsVYpeIxcKFIPIwz/6ZNYUsALu
CFIQOWfWtoZFL7lVhW5u0BYLigV3oC8QeNuuJpkV75tEyWSWxouBeBww8Vh1tqC5
6byH/uheSU7EcMD6DwD/rRbtnEM8eChsyk3ibQD4jcqXSq+NNPzqia65QBJfj3mm
0RuraxAn0C3OZm4Lo9YXI6xOIoLAEDJVzYBPhgAYPDJOr/7YuMtC0v33zT/wxTsn
ATK0TvQ4v3JW7rKzuz3/J+rv7CsdtGDL8KOIsoVPUmrmwNJbqyfv9w1OJGaiwE6S
+UjcX0mia0NTEJv18+HgfZLbRYOX8Cf49CTo1fGCbL1zML2li9X8qMqmgxrGtQdL
Ex3u7qStbD3zEeYjZfAjAiC4I53NYDh/McHtPc0kt28QfCfMecT0X+7Y+xxNJdIi
YT5yfu8P+JKKqA74u7TUPmRGgzojUwGwhjKUJV7VV6svoiNEfAQD4xe9Slf8BSJ3
TF0+lvS6oxiQx+BtarvMZRcRHFow1ZVE78Nq9IfbZ6V3z15Yvq4TQsE4QsB0nvks
n3zVZaHV5ULlCqs5EfFxjZYAw5lQy9fsmrwX3m6EgR4KxUSD3KuZiKO5Ba1eovA0
x7S50eaJ7HQRY3SEFh7z4yQUaegQEeodpnge936KrHmbmkcAeC3o/JaQ+ndhV38P
7omOchCpzJ8Rv9VsfoCOnYg9pa5O/hFqJJpiQR/BHibAK1aH2pzzCFAtu+y0PJpl
JUIk7SLwsxlmEvFon0RIaQhQrhBgAqPWzT6NnMYHS2CdPSGDZoe0nbsSp5lxobPh
fS2CGe5ychUfP2767b5VcT1qpKdzg1C8nlCS0rFGGA+MJqIlZBYEIMNoiSiFXoay
0D3tRcUa/4PPNUn6QcMcpkyQMVNyn2Q+STu+XjscPlPF/bBSoclW5WYogc8kZ0a5
xZm2AqTXtL5RXImHRsL/LSs33ZVv7dTeFqQxmKoKHQyM8S7VYJzEBTUf16FyCNO/
uR6DHpTnLEvlSkNU7Q/rpcl94BP6d+MQ1jcealm76aBKQMzBImarDAhx2x09wZ4F
JXqqxM/b1QWs23t5LzCC2bTGOXrV6IzsCVKGKFj2Ui5VDpWumJx+gXKcuIQH/pOf
dmsL8zYKaP4JPTtWhaXtag7twES/znrKsI44U5NNHg5ndkT4lT02W8tRW8n7g5H9
mH5DH5drdf4PjcDlpGV9g+3bihYop8x8EUtcUQuNnpHWtoy65r1GHIAH4FIuwuAD
bdQ2/yNJw4fVey7EDg3DT907EpamcGGcRmcs/RPgB3Rzd0iieqChqxNUk4wF0Xcy
RenBqdzQqCC6UeKznyu7nSaXAW2bCZ9fqfd+9b0FlodR2BWSCAa2ncTWVGIsAuHZ
puCzAkUXhucuyLJ0T9LddSNKdQQBr5TunQG1EjJAYPQZowJg4THd1Wp0Q2d1qJQ0
4ZmxJ2FGzf+547oDqpMjmsu0W0KYvqhSl9tc4mBGSb7xmgNr2DW1hVGf6U/lfzpb
CGrkZYJmAfsabRmCEPBrncXjYvoCXhDKeTqUF4qpR9JZUNjst5tGXU9b1y6QvhtQ
bEvB1Ac+Uu41P1U/yMpYtFAyXYL25c5VDndcbxQONgfbg9orzVemV9zYoX+sohzB
3RZCE07VaIsqn6bUTbNfKHaOOvx2qv+Ghw/JJU96DAXHiGSuVQACndCD9FElLAEn
GJjjUXhHbwMeQHH4jNAUDJj3evrcJYrlz1EnpbmnaE1JQo7KPTH32i2Mmyvc5hK8
eyhlEqimYjkQD2U5d06y8FqbIpj4yEX8SVrcfwJU6eJneAev3M8i3kyiIZEW+UNh
fttyQNVvozfa66Wx/MfMvA+WHX0sw2oI1FlClNBTPDySVoAlhAdi+aYZ5VEx3jzn
bgs58wDJrrm6o6P7jgXSty7bifBjhPE6p0B009s5yLpVOX3/nblL6zwi5FQXVrQr
vJEVu7ukauR05oQmBZ2DgN4HY6l5MedjttQk+18ZPA5xJvKx0a1lV56X3QycqGVC
ti+mp1D1JcaCA5HnGaZYQlouXrfz34NeVwINHa5Ui97FWIzCuPcRQLWPOEtYjk1y
FF8rNYn1sykqD/sUhFvA7zxezFI9uWOZBIL31iMKcVMiOGhcfOwdWMl+O2RUpFi5
aNEiK2X05YiWL+H2H0gPFBJ6FIKEkkS2mNlBPHHIdE1vcFRllbaN1TQlhR30gBrs
+Kwrzz4lEiMd6wsKpZlYu96Yeo6tUsdnkWYRuLr4NqurySliOdnVytUqfPWrDgQQ
QbvHRvWmVmPhmYcgVyJwucHHIeynt5/6SNgSfVUFVnwTwWxzyVgnRUuCvb8mlYkD
ctbZYqYMDhNfWeKcDwZCrxsnI++flNFzqFldanH9hDyH33GTrsEH/cEMQVRqu2l/
tDdQqVRFp3nligruvI21YRl9HN+VwYKkukgakCpcljpESjUonw9yblVAdhwfSfdL
nHIsRJd8Iys5a/xzytXX2+I4n/+eTPNl6MnJc7uIgYfxWWXidueFACIKB5C3aAoN
8bHYoDP0KczLmfjtjntQkgR7pIRLnstxN4StE7ahFuwGswAaCjz0TKR1sTcUSiBh
1R9nhMYRceEP0EHAjoP0X8pOFFrXSUWwMle6CRwE4b2BuWlnopwEm5x2GnyyT+u3
4yUnpETcYKuZyueut8awm8PDIuVDkucI8ImZRZcAM09oOcKoBGBTReB4XJuc2T8e
2XpUkL45of3YSEzESC2oKV8WZUduUVlZPLjs3pTedp9VjGly3Ytj3Guikex/P87L
HItxEPa4G+UtAP21HQ1BROXSLErxfspnBmEiIpQBB7MOEm/mOuToI4wYg6JJ36ag
nQ4RArhh18ffz/1n6INXEMngskqKJwZuxh0CJ3LenOjtoHD2c2Stpb7Bsb2pO5Xr
dMRLwmPpGFgQm1oTsKXagwnwuKSYPInIknXyJXamWyeasRWf5ZtIPcM70gCJ5rMs
+fpB0r7mKbCvLhLz9OaWkASRNwn994klme8m+NyzcrBw0sy2JZmeBi5boUa7hiYD
MRQYg4C5gBVUeksruL4r6p38x614TyQufibxnsGkGO4Vf6YbJd7akZyGsO2MV3qT
uZXsPJCDi+Y5iB8Cypx3gd3+GS9zfNZ531qXtXJAdwu4RM/zorCFEnqRJ0taxiCp
DUnf+riYwGufVfCmZnRpTzVGMzhoABn4BViobGY7RbecxW9Qw5bHwRvY+IAqKVLH
ywGmP+tpboIX6GMbY7BeXTQjv23ZSCS436RSIyGo86gQdd4yePlbh26/z4USKTn7
EVcEs0l1bBRasYMh+pd4or0I9HRI8urus2NWZ1qYbeqq84zR+SxoKdc7oN9MHlBl
X/FJsKU+WVbLRCY9TAhMtL0HCLqEeeON5PHYxpYCWAuAz25mitfpmlGnVUmdOXB5
8NBwdo+3xCvI6Pb7HeZTyvLeCYFOIZ/EVDdjlYNLmS3uPFvFMxZ4A2KdHfmOg+pH
/feZb8dTg2N01qzDQZl/Brh2nAFhvXRzjIWUoXBZzEH3e4yQe7xqcjJE83iyLxHx
hGGcF8dfi5wyw4ZioQ+zbwBez+ag32Ksoj1zHH2t8KYuU3oJH+8TTSmOiqnIZEHC
BK2BJ++jYqJyozuXc+++bhdYweng+LTy/88alsm2tJoVrzIk4xsH31kvmL0Xk9xK
amqzHLGUgVom8ZhEnpSmOnga0w59+G4/b1bAJnuzSyoN8yevYMXqdE3e/EElM/qk
UjO04IA5lZoUA0iGQ48K3yCzIOTFCJ+IAyVc4OeYNrLR/bInCHVX2FQmKjdeZ/uq
RaFCeJSXoC7UmvtYM69PvlM32KwDgKJAyxwA8goDOiXsyDvAcvoJRxhiZIQBO2f6
XFNdRb+rGYTqPcpiL+qQ9ibAIa2+MTKK3m20WQZl5ArgWKGj4ZVopYbnA0fkSMwO
Z6tPt4kVvmNBv8dSjg/EEUprxwI7FzTD4zQh3MHt3/0SpRXOYIPR9SaZYKKl/TnN
nj/L9tgCDnQ1wm1mboc5edQjKmGZ4RbTJweJRBZBahWafUrliKfaw4IvdLaGaDln
45s0+KIgVFwVwtdFOG8oQ1fAprZKY0fwIoQwkYA+BvrT0jJko9xLuulcwZYVEEjX
yj0Ol2xDFuXI8vh2aF2TcRP+T+ETuI1TMd1mdXKNgHuh1y6rF7eh0IbrZi564nOJ
gPqYRgKuZQ8X+CFDE4MS14GaOvInMO4zB6VSh9dFapp9+PiQ8kdgwqGiDtolNCoX
d+18wJbZBtTNEmeF4clG4FzE6N+8WMCXKV3Ki5hhBoyVNkLHoz1cEVufNi99iG9i
ZyzmXkivKoW6KO2diio6U8i/btqw8T6BhgKRPqfogRpbqPLOJtWhy/yryF3Cm6Kj
0Hi5m9vk7/yTN1ggclrJnw6E9uUKIQZvaJfPpZJap7CRT6Zp1mGzFhFh/g9yPlVa
AlVYBnO/CrCorfDM/ISr1/cN1A8iPOqryFaD4S4gt/k5fVuptwLoFQyjdY9Qq4bu
uH0iOby1BM66JLMAtv184izz2tuLcF2iWfBSg49/w5Zb29rlrfz4Iap69hfmcoOE
yxgKPNJTDEXkPcqSpK2RmDYMUjdmWLOGGsBI65+mR7QQZ6TJZ8MMl98bTkroOblJ
CJp3uj0U+w6yLS6WRYsF7BOBX21omH9wfbkfiWHK90XXGEaLQwtdWkJKmv61GY1I
W3p3K9h46QbfTc5xmRfoCGL6gx+RgzbZbUW2U3r0LqW9i6QMU0bFq3/XF8a/y+xE
NC6yyrQWwcbGHy+YuI9Gqa4jmmWo/vlmiA7ng+iwMvnWTZfdgX7/vLo2KQH/QH39
DoItmWb9tL5HsrX38hB5Ru6eBKaONxnxazb+Ke3kTCdG0UkDeYv4N5b+Q3SLDc8W
Ayz1gQnlH9Y76TUKBIQNJF/Scqhm24r58MPGghAIqnzDXEX+YooJLVrAaLKgUvaz
4sYXGMD5kJOztluxKrM9gJzZ0qQ6M50UBUQfUl902xVNequ4aXMqg1SXxspBCg2Z
60I4j/ZjMlanLs2a+ClRRGxJkk2py2RcxLXXIuaWHtB24u3nMm24Ss5DlVg5ZtWc
W9Hut3fHkb/XKU3PH1/G/JnVdctUQbPqQvsNPlSQitKns5NNXbAcRp0vgmV7uxSk
gTXTS85cd81GHJ+UNJC3ZkClVLps3tE/fYEnrW0/xlbCWWpDdaziCEHnr4FFO8ba
OcotItRALO5I46rEEzfTaqZOJsbz1U7k/oiPDwaGORzCFhM0wZxIaaTedLal1F8a
lzkGF6YICmooQjnXGR6vpN/W4zia8CUAY8lsAXKbsbDt1KisWtLC26QpsccT1N+v
HNipctwdqdwq763vNV89BIaQny43nCCD+E0rQ7Wbwh03Qwpn7lQC0wIHUiEZuhFg
moyUB4ybpENDrXy4PBGJYZ3YuLiVyYlF3GBt/ksWr1JOr5CFAJBCvTM4abc/rR+/
gbAQEgc9AomoqWMH9eozaCJ9ISBTV8+kc/LyMjcokVcEPX1Hmc7ki4zAS5h9QCr8
hwhesYfyhW2q1cr3bFb3wgBnAlJ2ZOIyjMUREZEUAM91G0GFLjx/hG6RQS6zE8pC
mhZ8RqIWILYbRqH7naw5WqtBATxnlzNUj6gKmbWwYAFxMUqrmxXFgcPyOoef9T7G
imFP9gWuIOeBrYXSWit8ZyD/Bio9jqSPvn+mvP3vDP3SSZd7ySgXUrrc46Gg3lXm
HHb06N0+5soB1S/xcydyvxQ9qh7FdGXQHTvxWXsSRjYPKmlHbYnKANh99p+JV6nm
NSAHKYjmDbxSL8vL+O7j80q2CRYT2c5NpC/ILl4WogEQu13ZAztBGNRVyBDU1ReI
+cdL0SSJ59L5ZXRH1mLd7mio8m5CQK+b/56UKWt2ZPgPmeoAQzQ6KKqPVKs9TZt7
AVgECQSV/j/7qn2Pi46JhcVj1ipppD2KWA65Q2BJJOXuD494OF8f1MmgAGdsqJ+a
Anw0qQNSYJBUN1MDfaJ4NbDxjDY/a2438ks7Nf1QAr5/IF/zvRIwkeKakc6YrQyx
PXZbkjWwSw46VWyVFbrbvGYuA8awrRx3EHG/jDeoiGnnBfAZQ59+PQDwVRV6SJid
Fb2NMVpAYALle0HDtVfugjNWi6yuIQOpD+pdAjSyRnsaDLQHVLceoDwYT7NShOZF
Tt8gN87h3XYUrRhkdhZEO1aoVDCRzNR1g3/Us52a99ALKuq6gts8ufxz0+hu1YEK
9T4ysGAlumocuehdMtWtegTrwMjDGtiyr9wRWLQ5db0rDjdMLtF9v0U6Hw5uQYoV
LgkDh4kaaszE+QiA2UZlFYcz02LFKCeDLKpxoNbTo+IyrqCN17t4rBURn8q31svB
5lgmWoEgFnaRnWowD4hVz554VRJU8lssiKzL/KTGslxdyQEeYoZOr28zx5PD35Fy
2rnaElfplfsMxoUsFPyuexZSNg0UiS5dLjvXFS8to+Ot8dAX6AGYxgpycLKO8nm2
YM2blr4tC5gaqRQgjoox6OtIkbolhz86ktmoeK/cpaEyr1bRl70XH7IQY35xPZcJ
Suh6U2jlAsLKUTsqSAy0HsxbE95hgL83t+3XhIYx0OuJKWUq6yJE8Sh6lNChiwwI
Nl9+5dVbW0BiQHLEnpwxvmmZCINwJh1rhg3KUK9ctbsQE1p1Xa6wLPt5WQD5/Mar
1wlePblC8qjFNgRD6771noWdYjwW7IDuAXysicDXctQX3YJHVrIfrBQ/lnLJrqxO
gRHqEayYatzBAyHvSADH1mqnHF6FiTh1jyyUh0eAQDeg7hjCe9zIk+dYD27+CouC
DkzPRpVKrv4c/q84CQkmjfWx0ZFBoBRUrYBVO4MI+yY5GDb78t83JZFBO5F3RNJ7
FMjQFMslhzd6qTGoi3bBZTrY3+zW59Lx/MpMTs3haYog7zYTDo/OdEwbczZTZhOn
i9d6hPK9o1frkYkuETGZ6AKw8yQGor7Qr7U/lZZ8d9T+BcFAorbFQt+UoLSZs1+L
3XJxyEZVWZFNYWK0PNwBwu5fS7nTrRntbVKSfDyPjrP0jaKAjgViyP1VxigNAw+k
I1eka8/274N0rglzOjk447xFirErJWDSs6Z/vXLMCLGOHjXOlBYe8JljcfRaQpdD
XOVVkonbiCCeKIxbmVt+ccL8EOe134cIBzRphLca5ysuOaoCkAfeZ0noDXavO+o+
gFZYvTyTQ/ykuUt7K86+yTHafN5ziLItF9NpiSSdXlG/2hpRcek4g/NbHK0jDWNK
h8pWaPYmjiLaSSwy+TEJ8vDM4zi0GAo5GfCxZLQK6pxFFqcOi/pQfzPfi8TuVBzY
AsSECASIZBNfDMqwfPuXIoAu6hWXFpZjWLHdQiyHCT7bMFHFHNpTv6+I3Oy8HO54
AaOIcFDFO0cB14J0VehKiQtL2Kp5YF0J2CgYlsP/ae10hwZ1TQFefra+kh0GhpB6
JMccSmtzN1rVk8Wu6GbnCkkAhiq6zDV6FOqg6KPAPPKmW1mOP1OrK9xkg/HmBB7i
Km7Iklzp2IZKENkIy77qli+S9fXMa7D9c+jVhJnB3MycJQvIpleYM3ZjhUNIrqsx
k33v0mWcpiOO+W+yOJbNHaelvOZzWrJ1kBzm1ns6/TdR3INqcd4FjX5x92kW/u0Q
xy8h7wQPHUORK8xDFRyMXiSH/75RAbiUtUhbS0VQfj4M8SPu+ry/VSimL4H5pL2t
uxOi5yC7gNPd1KsuI8v3hmDhjYoekXpjX4bUBzT8GiNC+g7fL5d8N7p4hAFDtLv6
gpWo3rN3BSNIh9juyYGMMwt33/Zq+TfyKlNGIP276SfnadqKYQqnaokFSYlKR/6l
W3W7Go/Taagh/cdGCKpnc6CVT/hylchhXbbSqJUbJnt41xrKuvsQlWCK+sw9kf9a
diE1+6IudjOFPDi0Ne7lcYESxx7ClDfOz9mxmDkekPHqCF3Ucrbxy058AJGDD73+
M97ccItH6A9m/rdRuy8GjmLg2zzlo5QkLBGZp5eRKTCxYD9Qz/T9QRaTp177Jo2H
MxUiUOn4g+Yn0iwSgJ5zhdDEv/qtb1xhNsx5QLAYXoDrjX2RojqoxEAkknm0XBBl
WtTJpv2mbq7/Rk0HWnfkFCg/SMkeCKPoC2Ute8hztge+InZaqxZYPgcmrwoOnTab
8qlAFj/mbJmIK2g7RV+lSXy9BOWes3n0sLlUeJjFKmqT4Z30g5YSGepH9l2APpoC
MehycrQVuxRar+Q/AoRJJOHQ71lHddtsSCMTVx7SO7HacDmrKahHm1YqH6c7mIyb
b83yFIrv0pmnuQqDqNZ513ovrr3KlG4BQKWeEmle5Rf9gritCEGPcRBUaq6FXUrA
TJk/shLnIvLnIwsFLBJ0mUHwA95X1cH+uLRCB8aYr+LEwObEbqm79TiYVOTBYj+2
SvZDWceJbhBSb5zTc7EVBpMo8kOKq8QUFqM8V238NrZD1qRfRCUsjnA546N4P7Sp
9oOG7a1yQXLF/8OAS9M/ov1FCh2iVBXtVP+GXRwLRaDOi9AsADqv/fgXr8kLoHUs
pyhcBAe3ILz8DA8gWk4+CeQ2KqWh2xAQJ1DIJ0cLP0lqQ1vI1iw+wmYe6V8gHs1C
ViajzKJnQ47x6/8Ahbt9aTfq+lUw/Ets4mgpCDeyZ1uqwOmUH5veQhO0XIc4nl9/
4t7z754xmX3RWhoucxAd66X+vmk3GkQX6r/4I1BOhS8Gs4LQkW7/jbkNMeghKgkD
iN2AuEcFE8NSkBNtgLipssn3H1DK+v7HfDVDr4OyOh5LH5N4yiPD9wftnvXhkyEi
tgnK6VwhqEeU37LD5+IKxFUze/+IzYkyYRclDdGi45MnOfi/7wKle9thbHklYSJP
w6oJY2eQCCEHm/I4BF92SwaAXtTqQEfSU6Z8YT+DANgHBo1XgojZ5E54B6jdOlGw
Z3QT3cfqWbGq0aIx5WUfTg5JQmB94kKAIu/mXy4DXatkfbKWA3N9aSJMsjeoRSRo
muTrJWg9zubFV22sCYYjEpjK/AFouSYIz5Gq66mG47stzC8SRebVNze9XMCUhMr5
1OK2cH4pWKjdD9MQ96TG1WXCtnCXqGxQpoI33vkVruRm8pqwehQQmSnKUkngBKY+
PGaRPIjSIN8hdQuj2mZyOnF3HMMH4uraQ4HvfwbUsJhVOlR6VirK4y96ZF6jcWq/
ziaN7nnvzUu4Ly/Jvwh8mo9DgJ7zlxOP7g2GrNH30aVDCTgeWN4dgnBGxFSJpG3N
fumBUAzQyKwbtWpkuSMabr34Ij6G4/CLeCoF6dzP/pa/IG/UciDSMtWPLoTjNOum
jm9z+ikPlpv4qh3BwzU2pvtP54MEleZI1TmXzYjVPhQmezdeAh5ZteFq/t2mgU3u
eoYMdHVTgQz4kftw4CrOUaEVHaCq/4TWNyrkAZGlbvlzXRvf0Pv2mcj/BjiM89nX
uSyPLpGqk8QN1ElN4yoYgtI/7M8DoMlOBZgc17mj8UtKEiKXgClYIINViKQlHYQI
P5r33tQmEdfehG/SCJnZvZ/nHllA7VQKA4xqoZDNKF8Fj5GPWUGd1CJpWat+M5qo
zQESCl7Sni5LOAGWGjjE9tq73URJUP4vFN0I5vaQSTvJ3B27fGJC2+0lFRLvl935
nlD6j7eUitYrwabDp70tSwgat1BMOT8lNZeik1WZVdYA2VXXTMYKYaAVgw2la0ui
NMI82OIKYZ6BRkIuSPpd+cZHm+lgkIypYlGj9Y5rNSBCtiilFqOa2LVm2GQ01Cqg
LpllGTeKiU0pFSRRw0j11sg9Pr1UcT/vnoe0jdO+qDmzLsl8EACzsT0X2KNAv1Ju
NJh1vMXR+gOw+Y0JeCyYkCL9WlaCrC0/jDtDf/ihWDDT8LM1l6wiWxEUFG0Fqw1W
ZNC78texMeCG9k1JebpQkCVqWHMvj9QoPbeh9vpXNjkCdd53+YNeICGavvSiRXH6
/Jnw66t0rOyJ2DwqkVTN9zoKYZK4Rm5jO1HtUQhDom7VJ/BlwwFrcY38bJglA4hr
82yXrYKAZKlazoTtpkZrn4ldznP74ial1+kA5BL7V9YHcGdCOCwZNE5mF52KSqez
qAoUg95TTxRdUcPuJDKwuenr1o9T7ojVfsTcZ3BVRvo50VOXVJ0g6TzADX96hc8z
tk9bdPCRobpF5x/G3liNgyTdKsok2QZkhYJGcHHHtkND3INgPefL0J8d7ehU3xut
6aeR/bdNWdQoMfvxxt+OyWodxt5/WCoD57oS5WBdinL7qmn3ivVoF3Y5RnnL+ekw
vp3H6rtQL58tlOkmIIyeQtoWxdUzDFSkat0/QItH99iKTQ56yiuDvmgxtx9cAO1s
iJRzVWqWxgXIeylKspZiVTzs/itPJzmgROnGOln3aVM6PWAawnce14WvggqtNHtJ
56X8Jps65/5DekYqZ3VLpAf/ZFL/D/Bd+cj0pW9ZZUEtTqGDYsvxV3Mgf1MgXU2l
4lf3Dwqfwt/xym4K/MFgke/NV03PPnBwMhMsTUi6WEPUCB9YYhYsnJlErxnB9BEj
yLYuZi4TSmODjNwPaO6qGhiCh6Dj8NczV0Bt+sjmHIWfUTnU9unw0a6RfhMwPELV
Bdo6ShF/IWiZfz78M0xhTxHJjMS/MzIGGNocPh6RHVKdctpvt9ujMP0uYKP0zIJY
o84FnqBjXs1NK4JSrEwj33Redz40+P85k/lUlnfGahPLN1gDfj4+AgWn+ZFShnYi
vdP+AWtIODQIWsAY00xmafpG5KAt+JP4p0SJHeDV9FX54mLWVXoFwNeoKYjYwfAW
Mrk4l07rW9uOYteWjxzQcdqA+NEJ2NnmrjdbNVzx3qzWwS7LTPS8jCvSlyRw3zkG
wzz1g6YVH6JHgtWHJvPoL+0ksg8iXzNcUov0VTA56aWmlk330tDaQEM8y6NA4pFq
+zwv4PGElgS6jfQl8CTIp9yoELWTChyUPcAEAh5lJJGD59f2fCs6av6V3XqexQOX
3bNSezWDK44OPs5bnUxq/j9KrqvtZf1e+OQ15FDBJljvX13cVtF7eY8dojXLpIah
GwSBK8Vj+pptr0ZHxEmKWpqIo4yeovX/K/sk+boyhSJ3doWq+g5RE6jLEbpp3tl9
+pMA96j9yn+LZebNPvdWautgCkYs5qEE6JDz+9dZdR1Y1HwX/0OlpIA8NH7+wTQS
9hOOyIVzDbvkLY23hiGuv3ncgdwkuUYClQtupJJL+wbyDpjppf8hLr1gQfyr/WZ2
w6tK9YnvVBRHvhpxtUTACAnrKwBqGuLa9kErMO0GAP/zVEfg7R0NbV1HAr+puQmX
rQHBrAk3qiOam7EfwbzxVY4Wqb95BuS4KUTxDSrMz4nRz09eBb8KSf7TW+2MR3LY
SKqnFpZQG0n3GJ0mVDaSHV3IlUKFq9AqBeb6BQy7q50yJA2WD8qq/xbVlHLUz5et
EXOUh3x5qPlgtPNrDOYz9AHMU3szsiEjGxRzE39mPoHEvowakYT/DpEC1dQRPodF
5ioZpVbmcwz/9hNGl/ETHzCEs8wEypOpr0hqj6rGEvQnTNdeRvJTziaZDf42gvZ4
Z9mn5N5sPyoVuf4qPgMFLFe23jAUxS1g+K78y5/XtY5k4o9aIqgi6qVqM6AOf0L6
THoyzUMYYyK3Wok4d4MtZNX6Hmu2AVKeQfZ+dT1Pw039WprpzwlLzTgHC8eVo5un
aWVMIO7ZkFuLbxkzUgBLmG3SrWqMD/vY+iRs5Sgh2U/9+OFmuMQLFflrh6h8Y64A
ihZE+gfvUqVWwBH5ugOSIKtYt7pzmKUBz0RIjjmmz8ZO6Rs+xBQba8VsBUh0ssNR
VgDF/SOTwQOnRYMzRf0wPu+pWT79zkJnnaLBN4CSmZ647y4m2wTlkotn56W9bn+i
tvREqXWZxqaTdpS2CfQHSD2c0eNXzuX4luoBVOwEde9s9SMpoi7/N5yV+32LeT7R
XBvzYCO9bnsQZTjvirXby2FM3KvWWyk7bYq/AZ80YpGf+29voGvzbvFIXTd4vvxE
PYmYKgB6tM7ZCpmiEBeyVnAz9VHC9L28icwRhQCwEg+nSxJcTv37Yl3zPhUNHXBP
49u4aVAyRAscYmmHceZsSxcdLSejxDeiV4Spp3ddQPUWhp/vFVj/D0Ro0zEiBw7U
FM3qYbolq5gSgOgm6RqpWowFrERE6yer/E30OzjmPM6NgMV2s6nGddxJgNhICRyt
KT9esV3GgsaBWHAnjsiEB2TDOLnLRzKgae9tIA8uWJYurc4s++vYZyfBm2VPWM+i
8qIn4oWXM4Yr0n3ZZujWBpIsz1/3AWPjiDcCj/J19Ft/Rh606ySTKTrk3zKJjChF
ykwjeIcQFukdtJH+C/GJzUBPR8XHYLuXj4vTnkx+DDLuwmUzBY3t3K5V3FDXlRU8
VSM9vtlyM+LQJyPIuRCQu56HumW0B7aYRlGlriISsFzg3m+l2mCAUiEi8HdK9738
kciU7dhKrP7KkuVKCzXlb5tKVAHu7E3fmdqXERavhdwxn+bTGbD00mLvnPjtsKNn
rinccpVWuM6QSnO4SmhQbow78155Cf8ieJAEWBYBhVEXY8X1VJQ8jVLvo6fOTBys
J1kYQas8JBuRE1GApqNiNTvSMa5UQcuXkeIeOODIyo0MhlyO9lBHAqx0X7API1QI
cmp/D1BhiES47sgUQwsG+3jUx2nttLj5gVgQUjBF81dGJD8Egax9RAfXSOcDNnc/
tkosU349lUp9n4IQz5l/B9YmoPNSl9ZGXFus44xKli1bWhkJ/ci5Tmu9ontKy6UA
fzzkAfXu7cn47qdVra2advpsJnVbygaScWTmf8imNUhz5Ve5mR7q8+CfuRnieSLW
tekp6NvTEZqQjKTmh4qH68zuM6xCgfTftZVZvRHywaHUoUJLfbIKQ9r662lgpCHY
0DwcI09QzRM8KjnpDjWHcutZMiARZOD867oDvMSpXQTSjObdqImbGTJND0I6tumL
7NIDHx4oxpluwAHPR0UDFJFTcsKT+GGgRC9/+TuguabBbTOOoWEJGbk8fIbgWCLg
mAM4Ypkvw1d/L6vxzK2mZg==
`pragma protect end_protected
