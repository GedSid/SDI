// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:39 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dSrRpOEW17RPjJg3F27wqTYjVvM8XV+shNcQnqsiDZi6qCx2aItQzNH4aWf2SsEy
DzlLIblzIMtZKL7Ty7sDiLjY70dxoCTxd3VWMGFQYHBsmbWdgNxUIBnIAcYl3eaN
csWj69f+ScUSVTiBHKVkDrtFKPCb0l6U3Q2Y6PGulwo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1760)
LQAU3FcUYzwIvzNW/z3lj8FYbqBOLNA9exQ5jvLCjXrmp4kw7L7GJL9bVRmP5U05
U9jsycddSZUonWk58VosiKJxdjvc8fZTwnsa+QC1AUGR7pzLw/EOtYijBpW/SM6x
YUHwCCOomTNKkjyqb9PPh/tXZ99vQjSiiXE6at0wzJHtFQfjAlkFnl66IVvR9U/v
5IoTRm5TFTjlAtzVabY6PLdDjCO0BOymsqQAR0qpzvbz7TcPu0QDK60xx8KEDHpj
ado/juRtaWOUk2Mvsf22dtY6LAppirneN0PHyHbc5N/mPQTQfRPujRo9eUQjNWLM
2tB5bY/oz7MueP4FEkb1osU0w5pTCYfifi/2LWdCpb2YNAiiSpdQY0nJr7ZbtqG7
dcrRMM5r4xuHwduTpB9wX5J4PJXcsKxoCWTgdEzsEPVJMj1JEtxVRqcCPmZJeKXG
4ox09366GVd3YiciloqbjUUc35ORoRXwiJAeB9p4IzknkBO2IODayPDU8cx79RNB
ZaH6vjXPS8Vjyg7anV7COUL04hYkobmSJgKQd3cph+7nDNM7Ogoc33SL/sBBw6wA
xB4kEmN7DsQmx8ByN08fi0sZhtSNpKu22Lhvscofd7AoqvFCt8jZ+zevH4ApM6wG
Tjj7bxkhdc73qHhJ9jHeIPiuUlybWZvxp8uR9eDb9h6/GfdtZ4PaYGU55G3fcvWX
zL9vkDqPn80IzPIY8WpWhSxh/1yJPYr7YwitgoS6griwlqENMLHfwDEB6gK3OuG3
YuzhKyvyu7bJoQuJdcSZ57Ghko2XGfPntlIgrWFBDJiH7b+h+DZiHabNfr5Tef+y
cpMgVtO+ytJKkrDb2cRbfalDAS3kc1hINM6pMg/U6u47JEzo/HbJSCMTznjeViGe
il8qMmKkm7VXAqRGlD4rqrIFpQ5UYr8bQNAX/Yz+aO3MOdu4lk9lDZGnlAa2FOqC
MwpA/LhBvMMp4wOCCdqsNir5XNDYN6cwHQYwAG7Do74NwGsfZ1PmC2OPqrilm8z6
N8JCvZz1vmKrHZAQeocuHH+3B5vOp1+2swk+9hn3mCBC2cN+EOpVK+d40BhX5MHV
qJkzCIxoeTlCNT6VtYf04tH4krhUTLORYt/YMojujAuEXTsuJE9HltRUjhKMEDeq
IBzhdnklZFP8axJEWmUyDG867iVf/slyQAVIPkYBg7sPnSBTrLO5dj3PHTXtoMog
YvI1le/oYGtvG+7+mD6/6ywtq8odwkox3/ZDKhq34T4zmS5GyuUn/Gojmx0rygQG
Nht8jTv5vqPOGv13aGnvo1AaMqYdXUudF6e7B4pwqS9rciIU9J9QzfpQi2w0hKHN
OrQOdVRUPtt55mBSH1a5ncpMpAtvWs490t6E3CDdT/1EXk0O66BS4T4cg2GZ0gmc
z7t8FH15fgO35gE/wE1raNwJybbyQ+Koi87rggRoHEpIRlHlSdUUg1dxZ8wWehRg
NSv6Eu61G1l2v8oP9BImf2dLN8axdmHSRz4j7UcNZJpzwqKGuxZCU3npTOt6ZiGA
+PcUmcKsjNwU7CHu1Kl42s8v3WE/fq/PBzXBtNmj/+og584Ac9GsbY1j2pHNZNtp
YkS+D3SmQWGYcdca+ZBjfVZzylp2njsMbO4zPI7g6dy2d/Kxf+Hkp39zM3XGU2I9
ZktoDhXOzdQ250JugtdM6md6weHCIIVIXGzqOsiw75NuuIk5y6xnIG9PYl7N1Z+F
2nBZZXF/oCrS8m34EHR8kjZBVsK5ZqNg8V72nny35+nSbKXzBUysksBb/Shf+Ql0
xYK+5ChSBLMCGLI1JTn+RRCUXatxRfPLIDWo+WAw5CpeeIWwuxhkyki+J5y3CsDd
Q0RdCVLE618BgN/vkCP0ASZqvcR/sNnoHgEf+r51Knq9M9ENsFRur6HOLbACJByj
MVntkSEf4EmUR1sAMoQ2hnnXjNU211b792YAIVf3xwiYo/cztkm6K8FAqr7g84ne
Wct0E5uE1t9HWB0ykD+8zjr8kqajwA1zqJ0S5d4jbnv/1S38HmV3ETIK71mdzqLT
MmeJyy7T8rX2kdpQCA5xu2kO7ZIMiW4J5wPAaltW/O/TVNAJP8OOaXnscIclBqWZ
OSYiws9bJPi5O+Ddl+ZMDaroyehUPnaoJt8JvrIu2OoKmWl+UmaHhIgnd70b0RrW
/tJYt/yhvHo4/jUN52ykQVsWGxszAF7MpDLbr8Jup2+K52ExPkJX8/mSABMMk1jZ
5c9ZLYC5z+WzP3Fig3OcIJmeGtH0FXKJqcS56uzMGvsor+W2UuSGlJo7l8MMs4HZ
LvWrD/Z37l/rVp5vnUAh0Qa76YDUNy5aF1A2QvAkl0I=
`pragma protect end_protected
