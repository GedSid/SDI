// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:39 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bgqpSNWeGNPiME+adT3c2qAkT+nMkUcZjev6QRuY1EHu4wUMIYPbLW+PT29bngNe
SkCh5CMd7wnEkrP8N5SFNAygSr9KpEBcv3gfRDp5TMDF/ayO0QQ1m3ra0vwxPfbl
UUNS2K6fMHMFe8l96O/P9Ae5NFvmsqTJdwJQdLupJHM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3296)
aKKg9K00iNBCuOjZKf68M5+OjIjK3MquyICOiLyL7LVbIlTaLrKwvCDNhFCIc6KB
u+T0MUe+KjrDY279Kj8v7xbwJR5hdv4OYOWjsUhI7luh3yb3HxWt053+CGcRLd+7
IOz45pNPDbx9hKwwT0ZcpWJX0EHxmHkRW0Qts7sRoEj0QCXvlg9zljgn/iWLJkQp
Nhi+yZwvP8l8QvyB4HfFZuznZ5O9ze9aNJiW6EFJeIV+U6BkpZZMz9pl48psjirP
1HWesrPkLsVgyyg7C9bLB7O6PqU9G/RKmFdEqKdcfWzQe2bTwk8rnxMuQVRhEFuN
GxJ25bBw31cSJIqq7sEgVLa325z7MO5hQZM1rB62vZfMdSPJ8xuf6aVtXgRAcBRv
WHG1dtjq06uoHeVv5ce1DbxHehel+RAGjRlarD4bQwD+aTmN2dvh+O56eIpSyld/
o2rMNFEd5HVIcjxDYv5Gg11QOMov49Sk9hOXp4xjJquVGSseMBbutavJIQBaFLZ/
LiWSuPWX+DAwi82rsO+jcBs2Tw5gE7DuZiQt8qBCy+Wvc7tWjpZpGHp/CbYkRw77
+lgB3rja/86jw5CRS8oMUtWFMlCZuc7L9+Ywa7hzRImXzMLB4UQbdu8pkTtkJtmf
SQss8P20PN5qCu1l0+BpUMTkqriUE5cgxQnQlV55b5Q/XRQAzT3QAxMXnvBziS6j
4feyrC945Cwg6s3gn/tzCOHCzcLzMeh24Ij93RaTjf7hS74CNhg3bEwi/SVcoY+5
gDEWkp/rjlWBcXILUxF+RSmpNQn6EmT1UXzPFmclGHCIedLnxDVCuqcHXmWkuTLv
qKjixWRoUDQNLJpuUXx8IFjZNXv8nc5DFvPCxSAqBZ8wPghnpR6rRkgMEgw9fbPx
sUFqfgRpe/0C59y/Iy9x7HrDeVlEbG6md+ow1R/phUTu2pkM063kO9ntZlCIyUDz
7U0DNYm1qiJIrjx/5gHzjb54J+OSZx8UBmta+Xr4tOtKh7YvkIOvYil+ScBS4Ru1
ieNnhpwWoAfL8dBTIOAchQEglvxMP00d1CAY3EQC5kBZC4BJrQVTHCqnA73PmOF9
1/WNChTKeWK+WL1vcQOe8RyXFjIlu+CdQgWx8CgAc2rKovXg4AU1VgtGp/wBICq7
mAVwLp2RT3JIU3v1fITBBnfJUoJ90p7O0SGitFH/wrUc8wcFiVMA7NOKNlkR0MDM
jBhVOJaPZOyH3CKhG04sLkomVbzbfJsC199K0qOHH15bpz3G2u1DZ28p0j+c82E1
IG7eM1I1x0ye9E1gnjQX5f8IpjNkNpdGGY1trGz6p8HknsHm9fFOu+hIj7G55a2+
yPKmtb8LlVNVtRgl0XBvn9XJZKHxyRFs6djgCE7O6701yXszThXsbnj59oKiGIef
E+j/aq6+XsO/BqDMtmO017zLx5miEPISWK2yf5rOpe4zznjkP1brL3v6aykIVuds
6T8YMbWgxQfPmYXtza6tLq8DpgoNZnOOHM2jbKjZniSw4OC3nZFVzaGMxlC43a6s
XYUTVeGszXNDVPAb2PZ5Tlh7MqQ5jUILJhLgO+LU43GUqTGcsyynr9Ev59GRAlRj
clfyJronJJqKEMuO4TyMeQPBb9at7WucH/UQP/zBj8HBK6FvsgooCYFnDyB+t1Pl
yytx+jHTpsQT+eycnCXMbWmugDZMfFdlPQu6O08SUuIKWAofHJrPMcae8mMjBI1J
mpK8JwLqLudC7x7AAauLOemtXy0zP7husxAHDbwFGkSDMIh2VUOssLMBNJ6ae1Z7
535rNnBhq5uwGAqjdueRlmEE64XFCybdIYrmAMgne2cNzsccMckeYAtatPXnbVPj
5HZd1FiBwNS0699mJ+vS47XUPygNaC2XF2OVyB4NE0tivbTFdtfFBuKzwoj0plhT
sJXbbkoat4vcQpk9KzAbmthY5vMu21wD+u3UDoXBxMegDEXqjYURvHRhLYao22V4
DXNjlbVO9RuRf35cZ+hlLwJuPbtfbSZFPvL8ay1tXyzKJAay3qFtCU92fmj7WbqB
s+7NaB6+GeZ7KdBEgULOUYmoyvfeHsDHUoKx/qRWFGqdhJgai3vRSnKtzWsTF9eB
02lDR3jlSoAheionoDlz6RB4kUDyNtkfrODp/uayih7j4tqfDVzeI8p1rIwv25j9
OGOTUYu8VyEC6JxvUel0EgdBJCcQSJ+n8FQ+D+HsSSJo/SDFCUzWeQwctpjJQ4HK
KlGPV+H4wTGkAYJMT3n6sxUcRwRu6M6n2AdwUKmYv/xlXTsUNaIMGjJzI0gzcAg4
NtwDsNx4utqIAiXoYTRj+gU6paGL6OgGr2h/dYtyV30iqeUkc1OCVRbKMW54tCvR
0uqzI8CsldpWsY2PT24QJrK80qHvXtQIHSdGkCQKWQ+wnD4dk5bbwH3GtsKgtCAJ
U1d/64La5nUZieeZR0TbYq64jdgwtnWlpJoSHg0ZW/wyY1Xt6s0Nv6GIJOo1uDtZ
d2JC8AGo+X4wVEx23iJ8Mr8U/qVJJ4Rcv8tIlDI0Q1px8fo3R9Ekm+kYwwC9jc6j
FYtNGZg0XxCPPknIPH/30huKjt20Zav+7F3f3c0xYJwP15u4TKSBWpTMFluG6bxh
1OPx5dyyrHxyJo2Ol/Hqj/5t6x5ps3SBVo9nQqNdw+ybFnbldUAQ1Yy8nexO+G2v
aoKB/zVnj7Uk5EyBfAYLxLoSuAH0jcGQDdMACg7rJlTpCBbfrOsAXKPsb6RuQyPA
RxsJjEMqyoXZXsoiMSf6flHggzbuGy66q7qw1DOo3xMquS2WWXJWWOibaJ4F8zSe
FRUtuRkdiqBl6R+aPeJZ7BhOilOEtgtQL5vGikc1STvHy9yEB0dUlATuH6BxoX8Q
POIZsVArVeJTjB3SCxv4uG8OmExEG+r+VZRlL0Jn+27CgVXT8+IjVPspJd9AKyVA
czUHyILgFk1jIj4VuFfdB2X8c14UqP1+NUtSZYGddEeCOHnq4DXTEGF5MGMW/F4+
pkm+ViFSYgYKhaWWwvx4GvLNPsOb8eVpVpNG8A2HUpJYfFHIjNbdtSnVi53sP0oz
uzAWgCx8F0q3YyebfCCdlxaAVqQHpv1n/oGSYJ3yva5GC4HDqfGwTxT3prheViXh
BtjcOCoWdCGdb4wC7Qfwvq0mNUohNujuzmpClUgO9q49SMjJSQPzVEaNuBCjWjXA
Q8fQtPW0Ub/pEa6EgwCfmsYv9sPnLq9103aPBx2R7RJ1sQXFBDhyJMVsGYw0oHO4
6t6JBdsQ4TsdId3c7pdIZajnA8BY0+XI6nI7tnXIA85fb3B0Dp+aE5P0CiWFpR4Z
514ItH+ZPLazimtMUzeu5BUJ5AUxeLDjXwyxZbRXdUiAhiwIeFaPRL9T19g1EiNT
Yslulrqtd4s5v1nDrcz/BkrKEzXoEwORS6Qn2IKBUFThvFdsmeaX/HBBV6MXheeE
m7Og8toikzijer2zPBqHXvuNge6TGrrj4FiR+q+L3x0J06m6kcsDFkXWIHsYA4Zg
sSZvYB59PzaTRFXdmuf+Q/CEpYMZe3gTandX/op8n3OWtbwmetGySf0ZnHq6lZ2J
lQCsnTiA75Gppbu7b8sLp1htVOCf2pC6EZt5TsIBhHsBCRsY9Ef79g677l8SqFtW
MHRT74sdIBD55HutCg6238TEXVd6YUM6KpXj7VP4Hekatcv9r3spout+O9lJbGQw
ohzbf1gF0IFYY0gBar9NMCkHuYuyftqihHO27ROQrpOkYJPL/7tQtpugZq984kp7
We0A26zCxYwSXSwjI09F7GKzogXDx+n3oE9A+e2yVaqrtcu54dtvK9lFblvds02r
T27SXxHM2Psf+T7v5c+iRgQLprFStt1vUiWzxjzzAIjW9Ztwommq8/QWa/PJKCc8
KRTEFN/Lx3VQ5zvZqg9GJImzluR6eZKZ+2//XA0tlHyXMcWahqfhABAEP2Rf9vBw
wVCYMYgLHtrfnrRTMDcWWVsuGbF/oFu3wGJFWmcpI+zeQGUPWnzxB+rtnzvTvFE5
4dXErkNcoetffrDDR+gcSG/EYU1RyuXoW2PspYvW/5t3y2fWLq2ooKyZu6AN/Mh1
9AYXpDJbnsRMq3aA/8IxQvvo+gyuEMEetpBZhH/0PEgFpULR+3EY/o+pN3cXGqs8
HeEqrHiMsancq4n9XX4H8I6W2L34bC1k4VtdSppCnw1Idq0k/SK+2L1LNL/tQVSY
0Q3g6GX1xC1zLTpdI+r1GfQkpVt8LCvV3M2twvfdRTCxnmbhhgv2BClMVQVAb0MJ
DIvKnw2AflOBKm0YpfqqJa4GMYDXJXiaFAl12MjbxfstpWoY99qfymmDQgF5JB8F
NUb5UQeXNWltESQ+xfmcMMSACsWpvuJ5PoZ9t+cdiK0=
`pragma protect end_protected
