// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:37 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fTSxT+ZXMr0puGyPpteIisvEuLNayI8YtUUnw5zcfK1zzSduBSjGE0HgIReg+/Pi
hVd8S1CLbWk1saXi3RnkyPquP7H83tsDoFJOZ6VN7vDmLPWsxD6v09l1DzRVfNJu
AoqER/4tmymE6405O3y/6TmyJ/V9KJUpFug3lcejnSg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 125472)
3HsVZouosI7c2xyHneBsGSfnPV+XvTfOhboh+e63wPlInIuyabtZIKWNbmk/KIDJ
tG2N16yjptIa2UONAZBcVJgp6kyfzXyKWzcFStFMrOSiWHv3GgwK3BFIocgTFMGX
nMnlXvqURTYIVm5lW7ZldkK8PEkPRep0YBYamI/YuImrpE9l+NxEhL1CyT3ieggb
0laKbRz5v7qjWABIVL5nNg4bCH8am+2x8RzSeBncW8KPYZPuO25jjCnnzW/WE/cl
16GEnGUat77jSfhIum8NcLFmtQLfGkicHGzW0gZp2FUZkNDUXbXIsEk0NFy/rhq3
n6tGvc8zm2jMc177Yuoo+O35Cy8jI/mAD5kRQETWWStGbsw8A61HtGxeBNJjDkmd
D7vsBdXyvU4Wfq235i6qaPALYz2Y9eh9Gjl6ClRg4XDe2I5YhaMdrrez0bnthXoS
shjOro/gNPRlUsOWVFnDozHad6vDeC8vb9cslT4sD2FJbeAz0wSXQcgVAzhoCDkZ
tdxMUXGqsnvALViWvjboZOJjjHgnAyx49/6cFq5dHQERmc7p1NOA2uaN+wfDT1JP
O+kdp9mk85dGVEINSDEEx8JkSammVd24a7LHHhLjMP98e4D/o9LJcYRRQOkUX05Z
moNe5Q7L3tBSQh1dCxBhDhYA1Tp8SqVGL1Qx79YocgweovmbMACH1FsjEpU7CSQO
HVMpXr3FNsRA+Aybw4nfeh4BnVg+JdCpVam7vlE4+sdaxF0Kx0HOHqQvRWDjI7W3
R6PyJZA4Htg6X0fr6WD1TSwJR7iwkct2Y2bJI6jUIj2/SVQEZyXIfn726xNxADYh
lRlOCYGdj/sYhexX5ocHB/lwzh8V2NOESKAkXrW9Hn3WhFDDxg/9SB90/p/zvlGH
xVLzf4c8GbMmb3RrNHQG5uAQUjV8SndUiuGKqxDleEu7YvFEUT+Q8Ky7lul042K9
xQDQA5/h1eEVGA4RB0NRYB7gj6MpRzZY47pf5dCZz07tiDxx7BkmOEBHNnPnuQFb
Z7gzeHeBpMp/NFQeaZi9szfVHQXEqE0yHxZ0LII5//pjNRV7uAxzQQyctrumMbjP
W4k+T4npiCdbzou54Hw2o5JtywQaOFm8JA92Mqnh1XWOAYoCHluUxwDEf38nNWgS
UyoYWTOzX2bp6FV5UD2ljqo2SRjgcIc3TrLPxsAmglLp1jvrHQEfdySzLbV3iUvg
CeG9UJoD/Q6KOBsfU/FPrhtwT6QC034obeIS/zRH55NRvDupSzfXveVhNoT+sS9M
0fA2b31TqyeA1Ay/rFdWFSrV6v/uvujuKMsvjBf0EQsz52DSjDq5xRpFKE8eZ5AZ
Tw29TvKbu3L6MDDsKPAXdlqsMJkdgUqxnzfteq2cROMzhmT40w/DMU0hjN+xk9X/
l22jmCUqBZ+ZdN2mgQJ21yvi/XKfgpVBqULPGxNoVEZ/H7piTbS9GWbFSGNTT8Xk
HMgnCzqv/cjWrIo+QnpWF7Mnqfu11Es+kEMZ0XcUZzVllEuYP4RdtZ8E0w+3nvZp
LbXWpsK+/jSLEcYrxl8aoCUfTvjhZarKqW5MaYCOMb9rvPoVL/gh6z8CsO+2G1Nv
Pn3HIBasJOsRdCbKqS/rCBWE6kXcil1+B0Mt78CUC3Z3908ujMkHY9u3cwp+Rep5
mHWHxt9jrTd75AnyftVqd45Wna2JCH2o36G5xsyZETEANtwEy6NLC/ucLRw7nnF5
4M1cRUX2O5l74BIVWKPRwDUDwZTWxGS/UhyYo4L85UqWF5ZtUoLC6qFdR5ukGCvE
8itTOmJ7HllyieMuAljYiOIUY+G9OGGYDT9NjTVZces3irqqEJWeBBItJ7L1LRQT
JR0R0RrQNrrDGlVpFe/VMpNhGEsQ0EVP3XoipzG9Npv6cZtz+MGvIAXfIQIvsfaK
gvwmt/s/zrQRGg74J62zfj39RSz5TXnxW3iZegX37ylwHeaAJQrjIFF1Qn/qerD4
sAOZP44oc6UKtuSi1CJ0W5zn8Ns5ZhImiuZC+8mP8p/3ocaUp98ZbZLlRckQVp1W
Z+MffvYJ/xAZ3V85nAC7AbH16eL+qynis7lqiZ2o2MtyUzrbe7uy34gTidWl1DgD
XxUOu/ZaoOREk09NSBhGU79++QuyoOwXyXUgw0QPVpXbx5FBqndAQdloCsLoF25B
3mW37gEUG/fRuw1q3LAbglDomwUrH8+uR6uBF97PonOaJZf6qTKDkfH7pop7oxPe
Mtu/d35ryXVjvTENlaqOQQOQww7zC1ilFYBtCeHJhc0AqluN1EDuzaban+fhCeBG
kJjeIAkPPJh/LuzRNUjYvV5LNcB957Ig3CM6TqeVhmmO5ihpNqNDtpg5G8kJa19X
7boFVnOPzMdr9yfYHL/vZesIkigdjyxnaYDmqOaKz0+LTC8OL7qm91zT6pYArRrn
w6M9hJsIJpmaDhQuYGd4lPlyAaYwmr+IbPxGDgwvdCKOriE/T0ZOTAguu8zhq8Ly
nCSvyn05VZwdpj1f8PA+nwPAU7TB7kxvh4cxEA0XafTX9tvEqYDedNH5S/V3vHvx
HLeryiOuvhPv9fL5CDt2fW0lFAFtCAziA1YoJ06XGKFPYmUG3ya6QJnElgKSN0Mn
2wOt18xmqEaJDZ8MjUR9+6cTyBvJunFOMUWPdwNpXcONKG2Qh+WX1XlYy8+B9kDY
AUzR4QvKTbqfs/rs2PqVECSv1iKTsYTZ4vJOsr8qpA9ToK7euJz4ZL5H+QzTzdYw
tEjcltMn7R5js0RFx8A8V08JCMpVmWyZXP8xvMs0xDHFaSD8o5Zp/Cii7rFRMDpg
oCG5eL47N+h44jDrHqcJSnc2nGxXfB/3fmNe4mmt0nay1ZvODMLLSLN4TYaie07o
1MYz9BT5fpcjYCaPjgU+UqdArWthlIU+RQDbe2+0K6OqLeYX+9ZlqW0ZFrjQDDhT
9OUvo2q7LFRo6Cs6Bg3rMVLynZbQP3HXQq8jYVbmnl/dUTnzLAUVqXxn21LKQH7Y
yVMfTVMt0pVnzbseO6jWnS3zhsoo26oHpFQ0iyY7QEiQYEgt+UUvD/oBBfyLxcli
IUmfMkQsvxTE36WxpxVC2v5rhu4hSem5JWTUi6uj6Xk+QR6x0voDMdXC0XYCRGQW
Ph0MFs/tJ0E7HR946/Wo/mztmb8w2zoXYhL0imPfBfM+175q7bMBmXKIyZyPMCuo
YAJpLYUBHsXdz1fQ8yfte6TbGah/qEhvGXm0/f/vZqYUOhuIdlNVaA7WIBPK5OgE
3pHF/NjChXvhFDsf2enlJFcrhfX7wUsun/Vk40QTyGEhBbPZcblwzazGl4wm3VFA
8cuRPk5aJBLVGAtA5TJGpcRwr3cWWVgBa9iiSn+Dt48KU+TXvncHnjul+xuIGsfm
hxs70vX6Tw8uBMnr0wTPFJa53iAUBSswFBKtN7vZ+gNTcYnQ7/SZThlTkUdBXLIO
gmRdzE1Lk7u/E8Xh3/EkRfi8wdH4TbAxSEMyvgmuIinlAmoNEGsP7rPSHpaqTwys
qi5xOz8s1+WB6YvF+GfSn56fAohlAq+6qOdxm1JdFAzpmye5rLyk+ammD4pFKLhE
KXoTYP851NPASl4JNf6CAtQ5d+Pw+kROBRqVk/tm2sbEynCSct04Xx1T5/JDrbEj
6dba7wYGav2mSCr/BXgsZAhJdRqKrM1nUgLiZu4yxrXHX+nnOX83SFZHGUi50Wq5
d/I0wwrmaXP2GBnn1cN1MtOe3RjOLTSAT2DtoOdLoG9yrTJG+7zh/YpM4AMyqVxM
bfHooSxNPx7CuoXhWCen8BuSRjGyoyqQIUEJjhaBq96pDt1LECi/QxVTomp+6d9J
DEa+qH+2XNUd95rjzOmbRJYnenp+cvJPS46/HqfweCNX+nCz0x9IGmejt6iJWWEf
mAk1eMQeTWYac6D58O5Ad0MOTOiTQuhwZstcKPsJTPT3l5N61bgJoi5koxH9OOEn
S8I324xvHV/CnKMHXQStuszZFq/s6dhdstFp6TYeWbTtCiLS7mfurPZCdqAS9haR
2nMPm7O9h+IvbZp2gSt4Y9Ue6ITREUS4E8xHGFgjQxCC+xRsiTYIb0Iq71aAvUst
krSuu8AmvpCGveAonLH2Nh0IVsC8MEXjT0xX05OYaA4xbZH7hFTd4csAaXXj9uDD
4Trl+SVitYXtOzEMQyfBe+QQ4B8MQqFCMOE6mYWb0D8kNoFErqzXPXR2JIWcx/ie
0F3pCfd/MJOQ5bhM7EDw4NwfKX5a4hb0q68FZbZrTUtCCmd59Y4jQLsclUHRyQCv
ssZ/RCp2VXzIdkd4naBl+ZH/hVCSpXq1yOK/FL3jNxSdwMbfCBlmFxdty7rC6p0O
JD1Tp5E/f/LDpM65U8kCpzB+msEAqM1r3CnEejFy/v5HPNzqKgFzmZVcOETNeQ9t
TqnxTmCRazIHlGyhSWT+jI/BHMxgf15hBAf7YCCjBj8pIgaR5ZugFHWYJfxCbKBL
AeL8VD5tMD8CuHhq/1MDVlRX5QjwVaKxN2eAK2NGzE2DmaNBB06cag+u/xGaS5t8
MiMAQm1PSPPFezJK18Lpj+lDRRRpekQhC22XvPV2naHh+gS/HfqKwsMfW+S6HfmR
wyHF1KiU+mQRqsshYtgpkpiMHkERelpR1vNK7rs+UqR5yVUfszw6ylNaSWoZikOX
PP/cqoEERZCeysRmxglltGncfOSreVNN/Y1bqqHhypdEPgghuAQT+Uo0ylpsn+pk
cQrb9Qc2wjNz23pgpUwWT55X1yHWELTrNd/AcKZ+tuiEw5jW4YK2eaAlXlURA6Dl
gq1VNw/pDd1flQRyavO9XdSDHOfaVfOFE+vfrvkT1+kNpbM/+hHuev8nDBZ/yM+8
kH4jhqKilYoqyvz/CRu9lXT0VaBdiqm3xYWPytyqXeSEoVlAGiQOAOFC8j1NmChf
ZEBLCFEVSSvNTc98Q+sRUkh4T5JlCOhFUb9vakGUb9DIG3eISpECmxY27I7wwoPP
pvrcMfTOSNfOR7VGehm7QZwGtsUR5/ZvU+XOmx8OuEdwk5DpeMe8Xrm+qeaeO1AJ
1F6dOHshf3CACWZr/NXhvSfUhX9gutO0b3kdgLKHgNXI6Bg6hwZPikRDpqAX1zvE
ZZAaQVzRIn9maG9qhbnisZeo0Xl5C7sScJSQBD64fuDq4yN3d0QnQIhxR2EL+rmj
qr1LUMs0HXcWEqH7VSy1OOtR6vN7Lo5MgTOrdZCQOr/MVE5FUNStVrFCKvtXo8Re
GOaH05JZneQljnda4DNZNWTpm/lsqXyC6yE/FA8iqRldz03wfNbj7CUwx+Scd0pd
YnQYAsK02NKnXBUA7bCHe5T1jjUaqQPdCz+w0WyaBI1MDzyPcEwjj6kC1wUDyfsP
f25QQ3YTSU0KBgEtqN95mcwSiLC3l8NZpIHcD22AyTkiK5tkfbCsX8IJokS13SKm
L+i+ujLkf1/kFeP5U+KjdKbfI4LDwZ8YDAaPCuXEy0FJc/LGToCnISG92HneJmUU
3vjY/1qz8uGDNqrlqsFqK4vh3lVBQUSakv43WNLBPBLNARWnQTom3tZDnNV8XnEc
UaI/Fy16+A2B7N/+IR0UmAPmpoCx/PIbf5sQk33tuX82HQxSGuGnvDe150jGztvl
COCeNpaF8yk5tzqR3JQtnlrOUHWrPWd/8rtJNZTv1Ai3SSF5NyOwgZdVaxK8+AYF
pW/nPSaPp/J7BGcuGzjk0B/s8cWIenTKC17pKxlS8bU+CQekN8s1P/13slua35zb
ueKbyijSiwrp4mhazLXuSXFL1bGpqF6QHMXR7RRPJYfd3+XOCGzyTlbFDGa0ZNJD
k331XfibhvnLL5KsKp499X3zttApHDZkb+7QCXqamkEQ++CnCkS/PtKQTuMd791N
qsuqtFxH7I7jdVMYBi7HMBxN3B8fgLLIC2TxupnWz9UBXZW8PmZ2gYhOQ54NMylJ
HnRYpyQb03AG0LV63v3hUVIA6GePHw5RVnV2cocXdB82+tbCMihJMgNc2qVB45TN
V0BgJl9aH4Eia4Gs1/LbIcFErzrnMVyVrKy5F32aOknUqogzTWRYwUwoaDolFCR6
sQjjOxQdrq6mJzzXYkdgk7FQLZfMMQy5Dj7j1OE0Ia2MYZ9zQvg3/TuVfLTWKB9M
SWutzn7X9TUuQx9ZMAYJn7bV8eEMesmMx5R4+CNDRITwV1JE3G8eR1JZ3mgX6dmp
dVlZTA0azMsUrQpSIP6bO9vwgn7Nb5W9+p0iA/+/MBDezsVy9sfLEW4NgxA13oaj
l6zJ7LsNpLz4AHOdklZjoB3/wZI33Ms9n6AY9/wVLuiJ8BHZWOqrC26BKQwAZDwE
pm026Kvbbi697Dz5zANxn0s4KRC8ZwBN/Qbum4r21McCC6CMHfTc8iYpEbd/vq1X
OA6jFBYI1OXyawzafpTm99TpYPW9dOQ9N7s8aZjSkVjhoYhfJBO3cXMKGRV1lu6h
D0540gp6814u2zlO3xRh6Ey68KjwYkCWUYj44sAyeUWNiQrJ/LANpBTTw8YNZrxq
TAhrWCXse8RsOUMJflt/zd/FAHAoaS2HtRHwgpwZw1E8fwPHT1AbIIQmCW0zFf8J
OeC+gq5fprtBKpFemQlbQhCvthPguKnnBvlm2T9VwGfj2CEQWGiW9LIgHxhYEoXS
EidgdmZEBt3PAWp81d2KiksB17ElXBgvH4Pyg+uPb4SWXzBNgUuykoghdvksYGl9
HDOtV1e8rzAA2x9dgqcuGKkRIucDXGzFjC1zztTP+BzMCmalVk0JfR0Te+VBLVam
BRNsbDwpb98bZlXdYc0ltldL/+YynWxwN6xS2OxVl1CjKwfNile0nmTwwniiuxBR
8LSIIMLxI89EX6Ui+wOcy+iEU9WhM8gcTtjhDXTVhOT9Ey7W8zt04WudbbCyqJwm
D3NmkNbt3qt8wBGqSCWgjxyMTv/P8vA2GKn6SxM1CiFf2Du+ICpDQ7cciLcyc0wq
s7Pz5XHlA7JYVVgzi7jveKwYOZmypyVnHZSTrjwllTRf3ZjIheMpfnPuddbCnPkQ
+7suYjXuXYx6hSwlIgXM/NBZJmhUu91T+ebLe1/tAJ6s+lWIltSbjvc00NuONBO0
0UmPfIj5nNSQT/u8fygXr66r7AH19lR5CgTohzKKe2nZtUTEOkA1NDHvbtqakkNB
rZMVMPpaQSPb3idyfljuJhsinhMhab6hqz2x6JyfnzAtBVv2HqKWPX14Y7Ux1WU1
NTZuQz6D7COjwz1AD8BnBlwz4aNBrPBsP43sy4uC4gUaIBLjaCRe6GLcFQdTYNL9
Nfya8WwmXAuoRjZ+CWq1Yyp8nIN4NZs1eOD89QkQuleIefse6OxRcC/fs7LgqDeg
DJzhaXlDOGw4VIK0OQvJio1oxPh6j6lwRGTU+Ytp+VcDNHYaSPkuSXqjwyJNYx3K
3SF2JuTC5g94elXdxfMhXt2oYvUrWsN1BK8/6iqb6hTpT22ncKzJTwHLxKxMkTAx
6K921IaShP6EvBhYMd6EvjoCurYcA1F47+NubATrm1W/8x9/nR+WBcYObzewGRTP
ww+xVj4CAQr4XrqvaMHMjxuhOBWJs81PU5CfDDTNMAY0zA0MRJneC24Yd6f150S+
LdGtYMNEABG4eKPpAs36hAwi0/vq9wMpyBxZJwEJbQsHDUGjpg03Fj9cab8wqM88
Qrn/59lhFbQY9+wWQBUUfFsUqMfye9gDGEu1PcGOKWF6IRfBYSdT5bI5CDuvo573
0xPTBe/So2X9EjGgPTNxYb27/zXFo9rhiY6AZiypE9aLkME3LzGKC9j5JQSauVst
jca5FpBKJSTivVDA6ECR8XjLhDUWHF4iOZQN0PujK0tXtO1n2SbNkfmBfez8mYWk
NQeazlGN6AtNZ+V8dqb07sITvl5Z8WmMNoMEBvQ2b0pP+K3OCE3tFdsWpN1mcn7A
0QClOVkFzd92T9Ajtktl9IXQdXw7NcB1iNBLSOcZtDyaJSX+0TFF1XO9ejgFDbdK
dz1TdqZJYPMNf4sQlYWK6ZwpAbg0O1job70Ohwqtt4YGbc5qy8T+h/ClQjSboauT
VlWHJ4azSbf/e6NZVBuyYOCUjWiswen78fF64mWoz+I0gtP2bO2wCZdYydsIO+k1
8Tt4iekCOMcsn4IY+dFl66ZetDPazZ/VYE2SlhS2WOr1u9Bo+cs+srwzMhqCRAKO
oMtSl1DecAN7iKgvuOS5Z1lYn/2Cuba7qMpFG1VygeAvaq1SDO/E8XxAlJ+yO4S8
qVbTxaK7SgLFfWcbkQ8+heqk7nxtkE9eHi0nTuIMZ1LiL4cxVBPQ5R/Ok4cm1nUG
9WBkoHDJwBfd7bE32r+0NvqwImyXL+piTQKSgWi32FNGK62PMmiZKLdctJeskAEB
ArwLEmVGDinczv5PUZ3KMXmGXkMkiWV9vLYY508iqws0ViE03Esqox24dEdK7Ggm
OlzDdCwPua3GTbaxGzWOqJ4XdTdPWaW+ON7Wctyyqi1UAr5lxYqVX+lRusyN4jr1
CU2IAgltiWUpK0lvU+b+CRzS4A43EGzQGNHBHYzw+w3TbeXcUpkjTUC7IaaDzrQc
hXTvJddi7sqMMzlG75b8GcUee5EGSRjJhfyIP6pZHdCWX3n0LUPRmPiwZO6DRNZ8
9xEwu7lAAJ7anL0tXHPfur9Cwnd90N67nPuEb+nROUdGj0tq8577SoLdLltOX2wF
a8AiGj2fv6/b18zOyhiUKfeutgqQnm36JF8oWstS30OzDkYLMxXjV1M5DI6rwpFF
xBjcwR2vSWt8nb69MCQ7JSg0Knv7hi1o2rSjIKsf3dRuMyXtJ6NaGLFemzq0d7B0
GgIfd9PoeeH9dIMm+8hzVdd6370Lb+IDcpmXTlRuz6TL6oYWXsINcjR6a6RHF1ac
GGlW+9Ub3aeIitBuWP5NyUfKiUGt66T5FOyTwR5Rt2/rRGMSS6+pLdDnH4/XDmyk
WN9sBquyCuZgO1FyymF718sIEy4McRWPzhJxBQa3OZe0foIn2hz+NzgKXSMSGK+x
fmV7Kx2DokVZUFrLn9DRnRDD4zV5IwCs8EVDj00R4e2efEOkCccsfK3X3NSOVjmN
4e+CTWvRdrkpJqrioZ5kFv9XUNfzYI66tfmLk9mr5uEORStQOIzycmR0pTz7UApO
TOmdCh09+0Z9Ns91SmRYfd+2cEiYnCfwuzA9L0hupJDS/p5R9RfRSHhiBlNFyRpH
cLp0R/QSN/aOrkNQHWutWPlyjGZ3SUzzxwjOEYdRWkvoqCkhp2IbthEA6ztlRDD2
bs5MV20f0fVwYuYnD73PSYsPNN0qMNxEOBZ3al5ZTNmfe5JWm+/v6MNAzY0YnTUL
L6wAbjpuOAJ6gtsJi/wqjxn3wzAOvimwsCFGsrmNcAbM8CnBvgAzFRgvzqx9IzTv
6uA6qV4cNJtAwTMbhUnEHTQ+boDzZmBhqqdEsDTasZQD8U5Iw26hwK82hX5qHNYf
BX6GIOA/d7RRuw5IbraNDuV3fAwf5xSdy2rEmBpUk4XB8y/+XsMdEzWeh7905cCG
RCPG/I3gfeq7mNMXbrucYn9ST/0i/sz2S8Vbs7x3qDHPq6rT7MuAkpyc2Gtm9Ifi
uhOF6M+xQdICOHkRJJcOQOZX9Ix55PXtwjfO1JW45ndYSL7W+zLC9ihS36u3D3zn
FpWPSdu9pJH4j99qY9qV6OshZVAMFPONoH4uqEDKv4zDQH9VgShLXOLxiA9LjSw2
hF0hT9+Fq2lzVw7HuTtiihyiB+jkVnAD6O4QYzszU/7+GxelNiEkgVXsUEYxGJDn
S7hWybUrzQG4nctA/GVR4HY0aMsMk/wEuI35FZUrPUu57FKPEv8PhcaFU/KR/oQ1
61zJt/DDXkZkTuB2CI6xiKzsKgMs67KRs+D8odH87Kx3viSXGnjIOlGJiFyC1EgQ
a2NKVEiC/nei9iUgooJ/et/QAkJvMuqP1lXyhuLP1wdEhu6wvExADHNIKjvh5Xmw
TJcpw0P3rDTiQeOu/mbfEpuOseRrpwh5hgwXN3SWA5/fWOqvcQMCyOYDLbTCmXim
wnMMy0o0rknXRVS4IK600us7VSqvB8EcrucOqIvm/o4aHcodngQyjPASEa0CtIbq
ZTuVZL5wwLLhIz01o6/TMuqPRW6sRsbH+tlR4762tQ3HrCtJ+j6W94CbHf8Co/O/
9Gt2Wf1lY0BEL8mc9mURJHkVTsQgIwTcwGWymFYaGFmQ9IvNx2T7bYd1F2Df0tBD
KRHF4r2keRQvxL8s+lF5XcPsUbR9HdCFX6pz2BiDuAdu4o/uoQ7T1kn+Qxhx8KqM
68KdM4AR7lYiDEbiN/4GqQk0FtJDkGpNHCRxQqNYRPWHb2A9fCtu0LJE0mHfhI1C
pYM9naxwdlwbmFigIsZQclFBmma2gvWQY6Cfr1aqY83jL/Z7QuA+ND8ltQvVBZND
HQ2s0V5xkxGxAIUuJM5TDqMsp7U4BtCzuzbpsJXmxm1aa1otjqhI21ogCXHpwrr0
r1jFFZD2a/eOoeHPX1XIgo3nOZ4GqmyDjr4UViFNpVyksOgFaFwqPWS2QkyJNdcB
+Na3UsIN47++jsDIuPGZXw1+vVXhPVioBG9UghEV1/Tt4r3hDgqz7nPhwrgAckc8
FOI8DTbIA/uxbecNalyEH0e4L+M9+zCL4GTBkyai3/wYuye5G4XnbOUCQ1qTu340
t5yZ7RqJUS++Et1CnUrbKjczHc4/ta08kuHKl3oVGjmntPN/CbBe1rA97slnizuo
ofgMfZonSrkLTQJB24xaBMtwvv8T570ALgFjhsnYZjOvYHwHf8q27WKrnewyCuWn
WqPBLVv3SK17S9FMm3C4RSkj7xkLD2Evsf3yehFdLZIJs9dDMmHSihfbcXv+sJCx
T//lsEJoUz+btXI/8hFCujhL8yJVcYbwUFiCjgjXZdJoNnhge3Bm94rbf2dFzHQu
XppebTgfXm6mniv+5csG6sHLcz4B5PTt+peaw0EVz9a3NTuWmuq1vw5s1v+g97cB
7FEkCgj4DMm9AMW4wFZ43VUMLh/v2VLqgXG/Xcoah1PhamZRvj8rqpkMTkI2QQAF
QjOuaX9bMYVg0GPP9ezO8prsVBxmlD4kdXjveo7FKufmOiqOVcG01h8+CaUb9Q2i
FMbt7wz7csRX9gBWajALPxCFYPh3Z+S9rqjQYqKyrVbtINz5f7ezQHRgoefSXcbv
j3fbV16a3gDhcx1Iah8NmrvPvdPXX3J6iSwWmRia7/qo2bp3b2aV0Frc8NjWLVkD
Fd8jGIRbbyrOkIzI35/yLbhWsmH+6g1rKTVH4Qom3w460ibBnEUF7ft1VdQIFirY
gjPpA67l19zxsqIZIijEp5d7/RertDnYZ3FvTpyjTe9Kkb/nhmySO22RbpcHzl/1
RalKn+7OWdPBV6HZk4u/IDlp4G+DBkYdZm/akk+GBogBIqqFpAGdjzwPfu0V/oEI
r+pP0UZMejof5VBua9/2YFk4Z4uQ+ROcCEU5p3KEVPz9rOR8g69smMeR9l62JCwS
pIRZvq8kQFZPPAn3Z7rrs2CMPJZGj9J/7Tz+Bg2T2y4UmNWLQuIrIUTMwTrUHPgo
PGM9IQscFeHp5oX8IqnES/t+wFcRP6OoSW18hBcLqTXlynbXj82u6aRxR2vfm7mA
uHpZRAHSpKAgH/oHQP9mI/2SvkYPCMXy2lsNMF85tAtgj73meZuxg71Gq67v7yUE
pQ3HU7CRQ5VUc1uPBYIdo6pOz2TSYOZKgsw+azwSTDUJpcVCIQ+0nk0iJQY8We15
gHssIOExt5Ew10sED7Q1rowz1Wd7QdUmNBYNhhYoJcEkskCl9XuYvX3Ha1bi/q17
7C1n5tblHhVAeQNnQBFDM2GrNcWbT4CyANNIL83bkchQkZmztc/4RiFpcpH5uRoW
cxffyprToirSJxoaYvWMMZXzi6dROTmzV6VIfAHr3Jsj0LwO+wsLfJsnC/VhE111
6Wo7sH1wAxPI1CwKcQSXZHOWsr13mXM5T97HBvkOoAfRiWM4PBWTECYFWzYP/k86
Yp//67Z/RPXN2Pau+MiYT7WZdP6M11dnzKra7dGwAIlBBGz/hi73m9acc0CRAQvh
oCci0TfjJ9zx2etkLGGNn/7LftGnRxoScPm5xaNwQNdi96gI3ow0gwincOU3sGE2
MzFBZv/t95lkH7Wt35sibAbEDUI27D/XYowG8jzLFI4CKBXATRQICJFRtjEfdfaT
fbm+WmisGiNivUHW9pogcBa/qiDywjdyRfJ4NHXWYMTTRPTrq2yHCsfyLid7w2O/
DZKn8/Rdk6/JM1BGNSr7vuX0PtksTYV/uDKliSH2fHEioUuq9CNZJEgVow7xwWUE
4gwoBLyUF/OXJtRdrDTkFo6OFrrxOKRJBjf2Q/5xjP4xf0ItrOHePrsZBtaEKMs7
5RD7VJfE66aSE5H1mIL/Hu5qDSjx22NgliqmgDa1ohXs0fCYiZoW/q3sRFWcnTMy
1DZHcuS4UU0U6MLTkH70bnkzTl9LVriCEJoxCNNbcM+oUkHRayKBW4tL9b8JdsUu
UtYFNUlASS6c7t4iL2cRVBBTWXBF3t81cRf3N3tkDr1iz3xpiCXU1AsRduCp6hGG
pm1cXRSZzzanLvHZfbFgs0p//2U338cp2L18KGTO+pZrixj6JW+CzYL9THCXBmtW
xzE0pxWEfUdq83dvWXWqIeGT1VIcBGefe9BCn7SRZxJW7CwkVICVkXL/1e5OUM6z
H1GE5kvy22Iqqh+3z85EXueLG7NJJL/XNgiREoCAz4Dk9BwBW1m/PLwP0mYsedjQ
bxFSY3aiHNDAwG0mlWYRsXwNf5vVgzORQE6TA10C6LDcQP7PFfde1eNY59qoFl9l
vc+zAEzx4NzVN4gkn84U9AtWQRyW4oqArU/TDn3ghwJiDhhvsJ07AyespAcauzYB
B61C44+7UM2LIVXJRJwClsw9aFwu65qZ91YGw9UiEfAjNc41/4ra5PhMDYd+FiSe
rsis34iSKtXY0e9lWMFcKd5TTqyyyWsKbGS+LSeu2vwKyP6lrE8MBKWrp0lXzimB
XtVehAcmMje8XfrourAyuzFyOZIfXG/iNdpoIC/VyqUmegj9WAunVNVQuJw4jYAl
uYQ40UEHjIcUiYbK1IRExK5ZPYpxrhSgJH7nO2Q7gvHTLAQYSbosss3KuqXU9MSL
Ne39O92e72DAPj7UHXcClTduizZmNNzba8fqahukXUVA4P0sA4DKcb5wnxzr5sMJ
tol8mEIK4+hZfXs9CaKwDfZovSsJ43oKa+THRYcJSwB0mR1PCdlS+mo0QwvsUJT7
26gkY5/8c4epJ7dnHYXynXhnZaDnHtAa9TPpO8cq7q0kczJ4rAeXoEKXECdD7wqE
iXNgU8sngq8A2F50k7bzmHiLyE3TMaLFCiAGHOBWNzz+ComSRke2jj5oNu0e8rl1
0XktMWaWtJg7QcCJHHOEul+gZH4z8z0k2kPoQvLtPcME1CGobnxxNylp3Atzw6oU
EjCMh/xpObrV7Omy9EUoRNf3LLx+vE6wiEtoVxVvLjrJH8ZWItsc0cF9IPLMgYMU
5Z0ota7Ukfp7DtxwmM8a57XsxKkgDA7v4SmkcuYipvabCJSqjihN7s78whtWFCHl
3MvaF2ONPbrqkqRmUVOoWAnYj7t7Wr8UUcuaA0poank7aFe2H+ZeJw9q1wWvmndf
PgNmBXiQYV9oIoooXRVd/a7FK4pE77nRDo8jIh7Hz3D2CAa9JDF3CFKdjcPGtILk
naCGfULTK9y+11+XRusl47fXhD0u/Gp0PYDR7N78IXF4cAclA9aX64PG1F/PYtyJ
ns1KQ+a+UApCxNfissqR0QDfolFkvSOyxMvb2XlPf7HtbL1N5W+QisdTyh/OvKFb
uoG/cP/dw6rqTXTahxu2Yd0FIfJtEz5eD1W76zDmClGsJDnt+2UCI5/JSKuvd14E
M6rvKbmb1SB/M/f248sHiQSOQnoMWWoecB2QXjAl3QL635VjNwqwUlHsGs6yIk38
/k89ZkwxYjx68LpRk8YbCSQsG24VUs2jO8EDfciTGh94Ift0KQMdlt/s9ApJISBG
hrk8MafRgg4FSkSEvKjFxJZ/CicFA2/y8GLoFrGCspx0psZ4FYYl7htepM/iw7Ks
5Zvzo1pDGJ0tRxdDrdwulq6gKiXhrNgBlgylL0P8adNA+84enTivcrt/TyTitWyJ
xuaWVwujU5bkGzlrsESY4p1YTh5MxUhbD5ZMAOyITceWB2VkoTV915Ap58P97v6i
7IwJ25qqZUr9+T5SKnSOqh6uUdHIzrZE0ZXSDdyc9sge0sqGTP5bTsqNLqo4If76
aOT/TWoChBBo3zM8T57+zobXamx8zUZZyf7z/oALuRx0qALRdTI3NWooGkRrWIJE
Vr+NcTg8iYM5QepoHCwb+DSONuJAzvga/+sB7Hz9Wr2E9ZxLWdr1rdjZFCJ0UUTA
/eMmFVPlD00DwDPb7EvsfAYzNpJlfJN6NZlE6cSEvrBoctR/Fv/BcAY5J1lxs2Ea
cPyQlaqQHFXGMK6IbF+8ihZ3ornmDPcIW1hBIQTIIZFPiACIJ6oL6MSSedDpT7RB
dColwpJNJZXbuhQKlacnt/Zb26eoQu8RUoWCfq2dRCQps8/UcIzUny47sEYH34Vp
qXcwVXB8UqLLg4zoB9hiLn4pQuquYAtclTd3WS8IWEK2TkVxdBBVCnIyB52oYUTN
mbxrRGzKxZd7PLjB7mSJo8tgb4xwhkmRLxLeZ7buzntMJ78Y63p2awKhUyCQoOgF
pp/M2GzSASFFRyNnBMBtGC+Kr0G3v8HIaf3QsuHwEw6/8dkKUYfF4bigOks4P4x0
sGFoDoGwqlOl8L3hNTlNfAaYBQbFYv+Jduly/oxWImpLpAh0k+H0XDQ450ZM6CSx
vLMNwSOrd9Qd/UuU8tCv4jKEZ5qjipKtDXt90So4RIGp826zxM51TF5N301rQIH7
Oq0kN+AXycNOD4vetZ2VCrKcKatKAEJntLVS6YyeuB2lWWhGF0uF61iulNHrIEnA
OoIHgW8Bw9tCZRs6ad2AY5DQAQWLcyCW2ovV/AYYLAikA19ArRQftaWR115NrgG4
MAPT0Enb/TZJZpzAhFYklDN7NtbSh4/K+dUB9haX1zYUjwNGyj/fMl0nOrmgqMKn
XTFVTUeJmZiqL1M9+C30rCvG0yWhWiJjoSuDgTEG0LIxa88KzBBDE+p7EQqQy3ZI
J7co/F4Qge8UN+LG2cmb2RLGWe35QVU4mMd4RGtdeIOflLnfToDLpi4iAJj/227I
W1ZD28mDjjMOYGl8o0MXmOVITIh+RAYJz8cgggmix7K/lD/psJ2AZAA2xMpbaGRh
SSvoylJpKXNEZ/MD0BO8fPSsx74ShV4jUP6iLvpVIjDFmir3JduIlEf3khJhHGgv
wTg0m0MT1Kkb8dx1/gIB5qeE+KdxMTNMkDZ8mKHjVSRxrguuDxoEPWmtnF6paTSn
BrAaNDRFDPgg0KPwXBP1hnsPa+NiHMoXboNgHZ3CZun7ulOX/ARK7Cw2zquJelVK
6CZH5Pdxhn2mmJmctZ3VDCdViAonhBDc1UfsdJWS4ejG4NcweyI6KnRm84nvETvi
zOclFgVkz1gXbYD/W2w0+jhUkbDlwoD9weFfi42aOh9GnThaiDUYR2V1ijO5SqFY
U6S6qxxFDL8kVw5556aAb5Abobf0OsK69gzlR3Edzl5+JcJpOhWsS4El7sKhZZYl
NjyMYlv7qTyJKi+nL5lXDPVjfsynXRwGWvzFCiPZd/+GHijJHzdg7cyOP7Cxv3EH
ZIo0t4sXjq/6uTYIORE9QSguYJnxAX0SACwMmYdIABlnLizPz3Rt066OGdCR7hAo
S1VkJgcomeUZyUOSULljg9pgytuxfe9HWE5IZh1oDW3n/QX34RxwnZ9YK0ABQ6Ew
lxs0tUlucRGtC7aHbq1BT7meV3ILurLH3Ic8t3HNB+lsyfsiIt8TliPC/R/+uY61
26hQSyXTZrEn4cI18J7bpAQ9HR01PfusHFhZG7nYuNE/cU6UKuJImZNSBNA0ptkb
31+xN8a/iLB/lCVPFWuAFd2cN8AYEf7oq9+1Tr7AbYdU+NzMZA5deD1RKsNpSKzQ
APnGR7c0di1l+ZA6xDAskzd9JSgeYRPl81fbcRSioo4h8yjW1Fz3SdJh7TSodFzQ
B9tO95E53WTbgfMl2dHNkT15MPOWzHZre+fTYPL1wScFwqmGgA76r+pXOv6dJGpb
Gyoh2pdyw2Sz27FOj9VJs/oKQx0hSEvhqgD2Sm+zDCROE2EmGxNfn+pIzuhd1OhG
zJ6fe0YFLDrVOT53eA4VFH+5R3mC7H57MmULodjznY/l2d39LqDTw9hPjY2EX+BE
6SgO24YwhWWn36IN/KYQavHsek2XFNu06v1dc7+mA8taDBcEWWkZY4xsXTwyTXAE
ZdzuyHSvIUeKOP/Dghnk74DiXRA36WEgdK+rzI3KTARKzg02dud+4oQg6YJCNP2S
M0IPIfogDO9xPTkewYWWf5VCM2b6ww1Qrpab331UVtAzDFfP4k+Xyckcj31RMq/e
hT/pX/JTP0vFguy2ODdsNsZZ6raM50zb7lg8B01d1pfBgzYkX9qXv5+qTnbJQhcU
na4HhFDy/h5um2yLzKzysT/NFygr+3WCBOmTapj6ONQybko7V+SokZjcPp+mCev+
DmTH4tCFavvzacuLgqLWVn1qYyKiA4m4rck0WTpLswBvsKpsGxijbOTZ6UQdFzgI
akfIZKy3t7GKUBVgj+YgkSBREabXkBrDQMjgvtbvMHvntbVBn1lTcJmRpz5VIEZf
yXRBJRn04o7lBL5Jh/N82hyNVENPjp53L+drwMfYS39VPkEuOnTXk3KbG2TmTrSP
SwbtplAoKLvXjX7mZba5A8O0vNXYK2RMZYWUtMnke6sHywkYc9laAMZ3SBEVO1S6
PI4lQcTuLwo8p6bkRHlUwGXTM+8sPzXpGFqdAbLWXe/4Itd2FTrmAbuvwKC41E2w
oBePqtBeoZA8KA1u7ghxIxAa8BqlPJilQlZEWDUWSmA7BGoZqCK3p1zPNUIQ6DAD
rm6v+bUPq6A37dUGLbeFZx0TmoI1+PPK/pHUokZd4qQhAnpBUYRS/8jtSpF/Sfkd
XLpzRby9t+cBglvYwNQnpLMy1MTmytv8uym20YvkUh79jbdeXZUQnlsXXkZOBS+f
+KTbaCy+3kQ+x4P9upzwCPdbPIat9MdIssnBnoCnOy9YC3DlXWBAbSAddzHm1Rku
DC/C8w/uS3o+fzCFOzcvaWXHRxHdpXiQYo7VqQujZJ+xEG9zxWLzEqBSh3zoflsb
f7kLKx4/tECrTl3IoUc5heK17AjbyAx8JAEobdZgZ2oKnD/+E4vAn4kq4Rzfyslb
ErHUFJkWFMwwxNTL9gi1/daUtBV4030hy2kjdelQFUhjTrX9LxaYwj1zN9g1tk26
ZnJqnCxhoVBwlYW3lFP2Ab7wajUVqvfyQzQclNzcdBEFg0ZYYzk5w1VDMdLtJiAi
bMdLU5Qzik69kQExUi8iv+wilP7QzykQbG2nHiccvwxfUJjFPdURxTytgARreBqV
7ZlFAwQ7/XmRG0g2ozfRs04MByoqu+NmfkccxMaLDfqEG3jeyFF25Xz19RxJG0z4
E/MVO2802g7JNXtj9nfyBGn2fOTQZhV/0hCwvtdjyXcj2YhQxFQGYVJnEC6YV8Mg
Gf7Clek5T8i84k2Yx50ZuhnEdBzFJcumItE5qUJI3wCJ9dKvr9oJ7Wf4YWm0v4y4
BFknT21VY8yZ6v1w/cnUkt8NPM8z7CEUcFuv6wYLG3AVP4ymynt9k4/14FLTreue
o9QFeKbxBq9rzPlezfB49RGofknI4QuyFKPxWVOKhwUiCmJNCbA1aYuPvFZ6MwTX
9fbhxgY3isYtEz43Mp9I9RtW+H3WpSo3a2t33tmmapPBcwWy0LDbHQ9oOllGwMo/
pLUCS7JKWfvuJmIJLwM2MNa2L2X5ku7bzqQ7sExo2X2eUl2U9GI71K9vBC/BVCzh
QYyq9hZqbYOiHxKz6oQrWNeCyd048F1AA1KYTxwSXGzKM+PfQSEnI2QokLbr06pV
PvohliuMQLyaKw+VdLqvuuzXNEOZtHG4lwP2DgWpyjOOVGzFrSbh5NR2N8mOGmCD
/4aQSKB2ojkfnePZFo53WoJL96GQ0CaGWLSVjgY5FeQ8EnyR0sFOrRoXGe654VCb
cGIgHwx1fuT+ckPGgaZxXzQZwIxw9vZsDQrdNaV7TjmTFSYx2cl3+skSN+QMtwLz
Ij6A3QjKUFcRya8B+YgxthP3/T5dhyOlktCRMpjkzO6tV5lt7p8hFDlmOSe2nre/
60SLIp7Cey8ywcXbKhJ5dd+tPtQLDBrXwOzOjisEHUSuWmyDAKoj4kUxlkCo0tUd
Z3yvrE5RWzrfJTvxfgsdg595NGnW8vLLSnIt3vKOxY4o7/RXTbTPnBJNgrwAsEj+
UTsqL1oIuSCPY3hRC96xM+iFHIVYLqYwfqxGMaodJu/fg9b9Wg3QYLPbZABHb4gb
eIh4CSEu5AzPfwlrQ32PaXZPFWmluP3AZS0VLYnCOaKH7WF5uVq7jfoI0uaDETBz
IdA2J2EDoUNEm4jdfgdcW8Ovws8D366TxhAS/thh1lHUcpZMiGLazUyThZVVgvh1
e8sXl+6SwngFSp+2mCumsktkNrbWQxTVql4uX6Yl7V/O4yLJvtwTLQFdMRtIQNM1
Ke8XRVfc2SnDiCnRfGWkVNtos88/oil39wJffcM8Ak2gz6O2vYA1w/7ftPzBIrep
TtT3rPuc0bacu4tRm658YgbHNEU+C+bmQkZ6NZ2SiCzCpHbeUz8R56s/JQ4wmItn
vw4D3jAonTX++9zNeyl0QNWhOrQRara5r04EUoOU1KZBzE0LRDsfMr0jLMc7ZBXF
bZs2s0yw3nRPzgRQEIEHWdlSDfePSoBv8RzMgxViiz7HAS3lOb17mr3dbJ8kz3JP
7wxoVzG1mgDB2naT+wrviP0yZx3DPXmex+7tJzXIk2A9FvobwIerWsaed3Sk1NuL
9J0hjghleWqGwkYbQHC4WaXtKIZUb6gN06rK32B5+y6MJ7AvqC2/IR9bRMXxzcWn
ZLGyQFB0tIHHs6z8Z+19H0QRvMAttliTuwrJP+1ZnHkATULruoAJDLmAvY02ZXex
tc+CdZRBbaVbbrMh63EPUb8aWlz0qRtE7AwYCU5/BfY+TsG360GzSy1153VabUEK
3WXaM18FLRsfDgnPp6CtqYx196PNFGELZYYay+buY2kTH+VC36umfA/nOzj4Z1NK
F+xHoI2P72QojQIDOkury5qL0vdWyKhEMt8U4T/8OQwv0z31HGimJMjRt8XINfj9
ed50teMx8xn2AxXTRx89jxLw0tu97YhOtW7UY00S7gwc2bV9H0adhYfOVsrgNWfJ
rbTWvW3l+RkyfAQNMXIqT6R+x9FuIYsW7ZzxGyQNxSmwWA4rrIVhwboKvLn16etB
gvOs8/c7mpM2y8AVJgxXT1BnEjE3N1O6HyOr/VSDuyYVkQYuF7CPDTg1J9wNdfzw
nM/apKRkH5uA9a0NFsN/xleZkuzOeMysEB/7dlI34PQm/TZGONWLPNS+YX7godfx
H4I1BfWzvYHTSXuHILbfLF2+9gx9m3nu5O7Vmu8SzVN7JA3LDL8yD4Yf8+4gwx5H
zBAAn4mg+I+/+elCDneznSH/pocRNZ4seSjXwf/IFWNZmikbuYNvf1Nj51OK+QbE
AmhN/oJheKnPbEjp1cBqVet7/YomN0gChipW9ETJXMgID+Gu5T1xSR6s3bw9s//Y
9D11M32d6gOoTdYkGHKmHAXmNueFkaqoHtdhRBbM/chHtlguvaJlmTPHG2cO2jjo
eeBTZFj713s01bSxSv0JweQuocQdEh1teRB/HITyr7IgruyYYFEexkr16WHLt5kp
YMPGUwA91Q7+l547UhqdVx4bucoGOKpl1HDnp7iVKJz/FFx8JAz8qUkTX4CKY3Ip
pwY2KcXpa3zkL6dT8jon1/Zmi6GAaMHPcuv3zzRq/zZGb3waNafFUlw5L9S4bE1i
3KdGh5YKzp3Svp+cenRqKX3E7RZRxl4vC42XF9ttjF6CYH5Gg8+ZKmi7TiJDb0Zy
jqQJ4ZO9aOChXB8HNODN31Xo30ieXg79Y7aMwLltI3st+UgrT6sIvPAhskRQFrV2
RMu8ntf7wQQ3XoLIsu+zrl+rw0ROcAs7sK5HWsfcgrAtkf6yy/dzeB9i4ummXUZb
78lcExmPc0JUzBPWduTrtjhOXzTfzMv+9ZquLHbZoynuiZZsQhS/fXLi88TKbz5Q
XqUkDnHtTmWuga0mnuOhhAFazUDoQ66H1rzShPqwQ0fbx0WjXn2QKCDV3p8zCL9U
tL6I5vHfYEyySbpcwckraiBDmYVAO7OgEUyJy7yqpyfxwLojoqvhb4dVCDKIQ2Oe
SYwyoav3thbCyiWRqRSrQB484KYhpNLJf+dkdYxQS6hd5q5YaWJqMBgMuGugf3hl
2s1VqvXU1obDEAx0Hqmmzt+5j1WG0ET7e2bGMTJ9Sdsak/beKYx33fZHrNtVrG6S
DhMLsMENC2fUEWGyUlYGvAIXrD1QGxYSmgwaXnrQqntzsU4SO8EM4W2G9mrJe0m8
hIlIA+SNcaCrgz2xDjk5lKMpSyably4/VJhWIW60DI1aqjC7vtD6Kyjp3kQLanL1
WJMRwu/zfCMpK56oVvK1yTGk1iIZNcfhbeAMoeqBDlqOFio6bInK5XOU9afst9em
CjkW0t2nORepHb9+qHx1sWDrDqBfxFv0/zCejUoFABKE7CCjvTQ1bNBivylCwWQ7
HXWBTWiKnOevE3I16nXivUsLNx6bEkRboAwWnpcuPlkjlNogKFa832y2oaik0Tzi
nFrLfQnXnxF3WUsEadeaDsePtZdmarPlTGaQ7daMyYoeksG/whKEoUgdM071OA/b
dVbvlUFd6m5BxGibNs+tPM4n5AB2JWMWpvRCzqzG43aiNB8ZcRm/Q7Jn03R3paGa
vjtcoCU8vDXeNcU+Sjcv0gWTusptfApe9Wu9Cjf+fvVUuZ7yZAX/Egm2MfX3bQdt
7KX+p8WJQeWDnWaNWcOpsTmZw2g3ZYvzISusfxifnnPv4aO8hI42DobCCgOuCd55
tBnw8QAZXHAKeVBvyTzUq2JTtP/lruMmtowDWhcYCW6hiZwUuuwFBQ0fItHt84ja
mxr3Bv6va1QgVaRgZsb8T0mDgMqc+qJcC+fzo4T/rkN7rnfKskDySOrNupyg6HdE
8BKvBSWG5DapFEyuSLlaRBv9uiMm4tlQZ+pTaqEx0GGtUzaIgeQAgP/ogDKEKGgM
ZqPGfqiAjft92HCwbdHMCHR8JgFnlJ+ZEX6q5NQ1of6+igh2JCC0k6R2+cx7hJLJ
wUyNJ8WBi4VZHeWhiQjHC/McKIUT7X05z8lZLJ6LktdVEQc7FVtvlm8Vr5FQQDmj
CxJaHAWTRcONnO6XOGACdCDIRy6HSUgDp6ZiY2ufqOZ9Oepywh2a/rGX/sMeFByu
yQjGjh1qF2BGckQUgD71oaeo45MnXJ8uufzRBmhPDp5nf3PVh9pqMBfp3yM++9D8
PR9sk7BsABG35Wee8l2AroFATsUwz94TbxDEdZ98QLoR1/NawrVqs1as+G+GaHaN
NqHj5ApDsimtDM26GVVIIoK0qm0T6ZC6AGS4HDCDs73VxsILuUIxa68bYO2ecQF6
K+Es4psz614+razJPThRfT//b2QP3xHZ9bptiwM8poUJsZ21d3w3EUxUfgZ8GUQM
NPyvMqNPA80bP8vZiOiBDxyZ2GFm7F8HUZQQp/uUGQpp50gCzmGTVmY5UmvH//QW
xRHMb11mI+u9ezcyMspblea+tFAnJ6S8ByTCU9uCb8wQye673G1o91SBDDVaD7Gq
RSRsVC235zE5v7v2nHLt8XAoeDh1QKib9XRzrzKQ4Oxz3T3eCSu1mzo2VSUkXfQq
bI/q89mun7aFurpkyYaDagBu63ztKVUx5hB1ue95HibqOtnsbFA8XOxTWXwVhZxb
ZmS6UET7bdOpMnqFs8KHEuBdCFzGH5Nudowbw/M5Q48rSv9bgcgzYpanLfMyok8G
kOOLuM30kEsBLWxUzbyNzIVtC+CN0AsNjwy/SB96yKXtVdI9WZhQpgTluK5110nu
j4k4YcBrDaJbTa5eVIp4m7c+aNxUIzS0mXkDm5ZDmiWxNgDI/OjK2VAKwt7gK7Rm
qwbjXdI5BiZgPnA9f+YIa3qSQKF+/ZtQIM4B8KWI33kZL3rIkiNPTD3hKbZiEaiq
5ufuPSpwdO+XCGrUQ8i8nZ1u7K0IfSHMmfjWOOlLmmjJsbd0h77hE/hszIec6QnH
qIJofqQJWgFWY1XYvnFDbUomafv5fZ8cjJLxo8lEMrAoUvWsNeXS86FdTaowfA9y
mhlWDzRXtJi92Ev9mV3NLPQC4Mxf/tCo/U1TN1paLfYvq18K7ObEm9rog3CnQxfP
KYJbdptk8RBjr708Z0J1yJpXKwMXZ6rkXhWM3FxW0OiYFT8DlU1lam4jcHes2iXf
jlDPZdLrtiVRFFE19F+hfQhZOeQW26/RbjCciPpit2w4kuLCVpLUvSH9/hMk1cl0
YMTmyiW40NtXpDcqp0egmhKv2OmW3hPte0/hujkGzxClvrj8vhnxdg78q9o6C9Pm
FwAZIutitrrnTkEbeBS85qDRO2jV8MMWnxX+NnxsciF6BIJj/g5sdRewY+iK7ryZ
2ooW7DQlDNr23b6IMrMTyJf+HHNcEfVDMc8Co+vUBs0wu/A7DG9cgnKHHjbSFALM
rYDlF+7GteXLtuqiOqLbJqB1rsSSrRGYUQQJ2e4tRX1V0Yo9wot46d5lPtV/d4kW
2pQpOwPTp3/ACyWXM8QTuW22fvGYYX1AsTAH0FiUNrhupIxgraP68p1cXhfiokh0
vh2jHS6cSgyEc0rlSde+uU/YA5YGltNcYXcSI8O8rrkR3iz/ypP0JtpcJcByDkfa
UQw3rTZZeGy3Ra/gYxT1Z3F6aprgpg4noH7hY101vuTXeDris3h4FAkBVVdwCrYj
SqAGnf55SsnLfkxjtHPLUwptqv3FEwIphFQ/LJj3IJz+uGJDOtl7v/uTq1zjqV8y
MEd8ynuSEcaVdQkJ29ppYnXyF7t2ts4AeJZSyiSWMIWFIRpN53RmQulPts13qFAm
TlIYNbRCvTXaAzVtcDKNB4HsVhUcmq4DiRallIkF44bUFslTDM1RcUUkcM7WokoJ
dlKArrF07lyN5tjHXdli0wJcSXLkFAVpsUa4vKb2VH0XPYp5at4/6rwEKPmF7NCH
9NpAHPD3xrTrgBrFSr+dWXWIUq3cgImLto+LIZE4l1xGy0p4wBTYdoWSr8QGkuqT
0cUxX3PHYKHc/0H1ZAvBk0Jz4EbcLJcv4rblci0Vd6imgB+wwcRXoEzyoLWvGDMH
Zkj8Hx+iROT0RIyHdGz4E6SxTeAM9+/XIvgRHZBDXJz/e8YXnCMJVXs+If1ux0W3
uNM35wis///Omkt3uddBl2ij3yzPzQZW/sdg6DqMqZGiZOhiPjJN+4TEoW4JVsGe
Y9aSmcKqElVzKOCs0oqfsKZGHzlrDm68+do1djKW3aLf5RD8pSJGCe+E7gL8WldO
kIeW1MMVW1zkIUw7INkM8FFjZwUMhLnmqyjlzkYPqZ7fMgnb8ITFw0pOUcLyxCTT
UAxGdgRFqFEWaYjBdrv3fk+qSzlUcuU/DaNV+Lhnu5cA2vDhGW87WOkXvY/fVq2/
mdWb8R77a9WKvqXiW89EovcEM0xGofjlMv/Vi33dn78UPeLAhnYqJ+oVpTTO4xmw
6Vh2XM4eE6Y0nyoq2E25Ha/u6TSqUXlg1ZkkrgVqT+pSwQvYIxWBPcTE0PgdntPj
KaCPM3BE9hoVL8mCi9jn8XJnQ4u4XC0THL2MRnKVus15aX78/uO6EusT9mAZFCwX
e09EdGhIueRkwEwURK5GsxAcCUKxqvs5FsUDFIZ6HKKs83RpOagr31B/fuLqmhea
oUpx0E22s33nGyr6UHvCOImD+TlMU78iQEe0GOeU7lNQSR3l1nMJNms48hbiIx5+
T28z9VBF8E0Zq6f9D9HYjK2hOZbFrUCrAuzL5FpWbcQcsMp1CC7o4GKdWbJrsCj5
jRlYgENIvspf8iZn+5LTl8V9Rmqh6zeJRonnPH5D4G9Vz63DftD/XxtJvb1GmgOo
pZl5xeG5hNPbyVhajParwX24iKSdxXs+Dfq0urUbk/9pc0vPIWVmIrSWUEH0bL8r
I6U3XCKFtk6Ocgz5ARaish5QA9DGkrDW1oBkT99CmeP+tZsyL6wyve5V/v6EM/X1
TCTkcEL6Eyw2cH6frETFw6+bC162RENaQ6pKGQlHli5KnO6vrtblrk4sf1RIMK2f
YF0UqD3pPrbZJ0b0piQEg0uFbVjMEePf+co/cJ8dTG4C5n7pOEC/ngkjJFiKvYwK
MYc/Ua9vfthkHKAlfH4EOP4XDvqBoIFlZvh9l9wn26kQvF6/kNVgEQCM4K7ox0I+
gDJ1AefKyVnsgdR4dYipGIH+wlpktM6pN1o2gJ5/OqKkxamFnowv/toVR3C9Bgrp
3s3/keJpojjeJ+Oze9+snDYU0ptK9IAa2u6BusSNvbn9LlNnQkzPHmW2AromiS+X
jQFccnVQRsIER/f3gVW4px4GQsbljE0fI+rWp6xbGtbRZjskHBwA9WfE7gOxtYmi
Y/gdWtZLY9ldFcvO/9HS/IvRxBiSk1lEQOVfw8Zz3LNE8aMk5QFRyZvZay9UlMl4
5FVr6lPyshDew94ZebrR5fpvEw1TfSFK+B1YKNDsqAB+wXFqEEiBxN4ksJimJvWR
Rb4cDizWFrpouK9m6cW0tCzt5xJ8m+6CGPtEY8tGzNZ6d+pi1P0YSx4KxJqMIFjT
Lnwek7PaGB6GLZj6cmdEj7FXP4Vi8PHR0os+/nWGPY2AULC7m50EHTHG/stiar0g
f5RCokPvUjVR2QsHzHY4HSB6KWPi1b67kJOfXYy5MwJA6KgubKr9yjxfiQ0oq7Y+
lwR+60qEUhtlKHA6HKFAhQ+FEFA7tTPyY8QD7OuXEgJoTeoRXOgv8jLGyRKFgs4X
x7FUn9qgy7gUPBjaX6FFOzRFwSlMjheob2DRrOPI74Q1wLvTgFU94QeYQ18emLJI
qKCvlB4NRcHtOEWqFdD2Ioe9u+kgYqfd41Oh+nOnvQcSOkpcAtSjUrYqyNHQpAxe
SCyJUM0aAJEpFFM0k2v13ByR0A9khwLllynXS8smhK+oZTi4ar7K2vbgO+kpPU0w
GkjKa1oZLKQHUrrGz6rqwiWH9G73lC5g31h+Haorrdufbzj0VOWrbTxHtkzGHNto
D/Vc0GuEBBe+uiyKh8nExckdePicIhY4pq8XNy4ELCwRck5tTQydS2bR7QB+OdwI
qaRS8OmSf2RSA/ZdmMdrh9WV5FDAO09ZbGewDcgfSU2DuI1AsoKveoy4Se39oE2W
uNtIwIgIt1719udJpcD9cDku9u5K5LTWXhn14M0xr2+L9+G/X6Hsu2Vl2w/QjdZl
G4Rbw8ECtxuxIdh0fqsGYG1pZ7bMpOT0Jge375On2FRJ1RQnBKqwq2vRTDXNR93s
q/gIDqyLQk5EvUcTOkZRpTCUY8tk7trjY+55/IZO7kPKX0BqT+kXvPptGbIlKZXl
Ae4R1agAdq/uGnb64df1dZbzAxzP/ZSCLylhAw9118vR2kcBXyEeLXxaY2F56Drb
8VKWugP3V5Isf6vHN5kjSrqMBkHRRsPbWiWJgGdfCF/n6Ip/GdVkeH/v+GtsVaSU
Pb2Z7ZYqWgfiZvu0OmJGzXdfas+BR/oTGY+SpqkLfTeKOpVupbpguaHId8me0jDK
fYIbGFjvd0qK+5R8N8CmSDpy9718EaKtrrtD/IXLRtNvxMXqO+kC+balqVvIgHs1
FyTZx6nxJnZnUIfLbUjUMlpQkXH0Xx2refyySDKNCrQYvkQZ/Nipwmc6ftAj2yu2
iivQk42HTIwqLYfil0Dmp3MNaMAlrz42OVgWvQlEkWAIRBGb0gjZf9AUlS8nqf0P
v4ZQk3S05jpBcfl0EgChXe3BjUICKVzjWbB+VDpccm9u5C1jVEO4hF31+0yknPlw
iOq+2xtqo2dwgHJ6gjI6tvXxTlGTZMck198crq2ivhEDcK9YTwGZ1LTt0Edzqdlt
++2yqc+uq8C+RJ7mGZ2RyiK1uZ84cUoDmmtT/gR38C1ek7zjcowkDVoKa+kQZYFc
h+OBaliNZe5dHkg2sf4YmYLmCGJ6jOYCBuwBymhEN5EwRKx09tzKy6SLVv783HqK
F/QW0Q9zO+xlWW4uwXsbTEMd+VVW4+5GQ2wwfLvvtUIMo7n7AvG1rQ6DNFJxWR27
N5AByikLzzlTkdPrCgLFCVjg9prLLYr0WgkKB/ARnjahKLmzB2VSHX/iZQ2lsiGI
dW6dShxcOo9CkclYW4oBFhWGPOyhk1c1+HHYb/vq9pA+KVff4/t7s/2prpDtPx7G
QFdOehtn6xQRbo5sWlHQLWED+kdF7aw3lB7r54w07+CtQNYgW/PHVBY5wmN/2GpZ
He6le+/4RcWmQjw+msakkbabK4nkwShTOO7kgOIDWtDOQlVU19GVU0+ZuZe5t9tt
xhEnj6nf8GdFgWamZoR2TZw1bWiRXpyzYLnBzHaVBx8+kbBy9zrUE95tv7ZbYbss
xlxqjhFECTNdNGD2NGkReQ/fNxWz3CWWbNj5pSP694hati4M4F1o/MQUbS9Nc8OH
wqTBYcOndkwtqqu64d7aiBsZ1liNKwcsfrWAg2On2B4VFulG9V5BvfvYDBw4D2kz
2CVVv1HghX/iY/OyKS+S6Eddjj6tFsVKfUrdE/ATBmkp3VllyYgN/Yx8bcUPRWPW
Zly4W5ny6iK0/P8ENM4HcmGJMsUaCpOJWap4Wkx6SUSSJl4SMgb9OSenMa5gNf5o
+0pgNOjdEsUentHmDH89ouBfDHj+7l8LfCluhaWv7TsN0CDMf4E16GWa5dPYRWxz
wowvKG6sB4As+pxwhRpwp05iHcbTDiH4DVfsNZJ/yzW+5aCl0VNFZbHqU98ZbsV5
8h8/MUkHFhfTa1OfJFivMLp4QisJhWaIa7QBhbSJtRr57MkE4kqB/p2cRg9/x7mx
Tu/9UUlkVu9f6Yv99+8c/+0eQFHDHjHyS00FaEgz8PSFe08bIPneZgBqyT0UAGF6
xHbUpTqX35F4IG6rJDzHY6t8FCjeKqHz+MSSHMtW5vksTX6iSGJBCivIohhVGpui
RvwT+tci0VlvyDHrnyTSup9wcdTNjWH6eXyN27bai1MH/pKvXOrb+FoVfgbXWYYq
wlaVXKxRqsoD+FVTciqvUQRWRLZ7jv1Ls67DGuKDYepUWie289tznAMXExNVuy+4
PTTcC3TO/rEPRbKSwD3gHgjLcixrzaq9vDmQHVX1ek4680OVb95yWzVZ70tvDJiE
yWrcrr6+pMLWS4d3YDBuGmugM+ERbgFITa0NJBDy5gVxty8gbIoXQHRc1FaamYTs
SVmPMo664CDfM/EEeIZVP8ZkoQFG4DiSaA2PuN6l2EOdQgBaiuPDYSzil+RbvL9X
MYyn6oo1FrV1spVKo5RbaA1pvVJJoWlFAK2GBvVyfCs6T6/bAGUEHJcEHiWTG0UA
+uwhWnKHRQ6gUFjrxLQ+TiEQ3fbuI3PFLSiD/NGFu6RPTQQKc/7GhjE4/hLMIkjp
BeMPhfxxncsoO/bpZdDk4VF8tr3QAim5+dggRHh2H9XAud2x2cuKu9ahLiHgOvWM
EdBZIFLkza+pGV/dSEzIS0YAqO28nuGCplApRCFrVqRBy7RSpYPz+ik2LfjcfAJF
0HuuYHCPM04AVeR/KxILvUDLAFnYRiwp4PJMq1nq8P4fBGKjvlYcpPPCI+ZxXml7
6W2Uy5nEd+NP7bjBte1q6o9jiJyfi5LjDt0z6076P8+zJ+CIt5D1YSRzy7gEwKdT
mlTarMectwMOD7yk2EUM13jQnne/eq4gh8tNMfsnC2KhQwh8a/fXtW8Aq+nt4v6Z
qcihRRlEtxpsYZcajSRDakgqTZmPCO3jKVGEFTOfFepL03ydVpjzJ/yuSQlEIicE
aEHed+KvF3UUZBra/fngIKWCWyJB2LCZZeBJRYfFRMfD37SY0t0Mzg3RPka+jeLV
wNTI8IXHPYATIIVB6eY9etS0v/XB20As/lY16djGw6S7hz36TCPS3VJnqP6wc/Ov
vsus8+hVmk8SlGJK8Wsy7pY4YYgOBpaingsF3OxxpBZXsdB8FeyFxEPZCFkKhTBL
g3d92Zu2HVJpME+21SUEKqP2XvvjtKbDxHCq6AMWWiew6v2BKiC0uqJ+md8Kx3kE
kYeRnQrWQ4HbupJBBHjH6pgGydlWxtL/DNDLESuVf5j7bohqaYx37IZxb0cFkoeI
YSq2kweaHLjz8OPTInA7jfUKsEQEYRlMUCfbaRIBH1PLB7WrxEVPRrQ8is/xlwrS
9H/dHxw+jOj9F/BiF2ceDs/Wv/Zn4BVLlGM2tsKgLTmsD6ko5q6ZKIsbcODHKAFK
tLzLXZC6cVjqpWMsKSFToSzTCott9gbz/9ejtmc7DsW87Esrk013Sk5Gr2ionybM
oILHnqs5owDk1qA3RhfZzEFVOyNBmE4TT4bP2WIhfG5GMTYy93XYM9cbfJU6PZQ/
JIOptLRY0iXKLnTyIjdWbgKTz8t3KQIez2LCR8Xsc4UQzBdPGUy1s9xHnlBS6OVo
x+C3QoulZEejPp6sxW/Q+BmjpWD3P/S1FPSkJpS/enfxnjrelDuDWDueQBSVLyPg
L7SY3/ofyjxaodZhRUJPpLzKs82YIqFY22+dznngy8Uxjrt1NxtZrswWe2brpJ0U
Clax5FKwpV7RGRZQMJJpejg5Cz6RWFsdBLCyQPilydNdfDNeR3kzFzkTxcqhE2UC
OwQ49W+cDAPt0RZNojKXTxhx9PTJBHJVnsEgslZ2RURShh5WeJ/0v1AAxkCYg0OF
vYFX7dSNmf3haq0yrOH9uGGNZadZkR79/nN5mkIN/wPWBXc5xHQ7NR4xxfP5/yi0
C5xEGB07fVsG8tSyMkCAX4+EpA4qvaKq/Fv7IN1Eyq2BIxFSi+LN6VYwJOHdwW5z
BCJrOeZADZKIq/qtRCJ2VjBudsQyMeL7bDcr/b5PdA4ie4A2gvoLhPyxwjx/+P3S
dUhZ++vmcPvTMw7GDQDZQgq4SC5/XEyyX8wQKltMQWG95kHwDs/Jm1JU2idqHwM6
QgyPK1vFWFjUXe6yfmK1g57N+4Bxi3pv+TwS+jMu++QOycqF3uzvKagTXw99GBsw
6s7C5ycUhd4GDk1zR2x1wE1dYHWtZZIUD4qctBroppQgcWx+iEFBrmIyF/hSD8dZ
f/5l+D6y1Da46SOKM3FVkZUXHVlVqAHBNsxM4MEdYZgQofC+UPdUarfwskNN92da
XhokHpSjtEt/qgTfHU2hk1X7Whalh8i1Lq5Ma1fSBJ5aMtVVosKymiPAP3OqgKzL
4wldGkdAtiFa429SZGG5ZphNQ7wtl8Xwoe0YmsxCxFTJ24ePZEYJGylSvSgC60o4
+jr7240BIXlLlSWNTSjC35ICqe3KGx6TcHfSv2nrMHFbLV7P26mXXhystO3x1AzN
Thii3WBc5LXZxzg50LU42pqtyTcjYlv2wS0HqU/SxO7mwmNpEm87l6hH9OyVA7io
y9UMWQtEA7UHiDRYUEN33T2KAt2num26H2AAxPzScFl7bzqkZ0wUY7hkC2gpVJUW
lb+IcpNu0/UjxUiDSgGdJCcgkgfQc6D1uA/v9dIJdsjkwEDn2LcBCZqCgfqlzFZE
GVjhsxJaNSqQjgK/7HJescxouSBqYDTTg34RpZKi8jctMnYg4KVkiKiICCQQFLpy
tTC8Yr0baWWBNFYEaYHRwCL02W7J5+YHs6ha4v6+SHDVuQdKoA3rYjGYWlRdxGOU
Zll0KuPvXlJygH/Uo9tzT5hZUQDg/9sAdMTwri1OfsNmxs1vG2TZyOGMDHwoQeal
5lFG1Czh2Q2ICIHBFQgpuWUViPPmTTQ/eUJ4x2EW0Oj64Te0w8qzZyDb1mFOeXK0
jVPPSsa0qUhdFAvxfP8Vub/oFflStU3UwXf9/SRbA4Gt7c5zr6ZImGfBxzcDhTI5
o+N1Qojg7l7/xH0+fnc5VAdBrSABebLQ1oPlLxqPIYJZiSaBWPBIoHYL/B2Ef5g4
9iJ0s2UF00JylycOzPvBghIF+Zb44zPEzwf5ImNdjK2g1TKdXfx0p8rKj9jtfPgh
qzM8PFA+AQRNN0jKW+PNpE/cLx4SpXiZdTCJEfU7+M85cA5VikVlPXvgLU4jPoEI
xBJaUvYkBoGqDhzGEaE9/upMG9S+VC9CKVMibJq5vPPGFyqwd7TM4fj2Zcir/kbA
zIh+igmBFKuS+ojIkvtoZ0KcqSzu/jAkkxqt4hNayDqX85LfbbSl1bUbl/vOSijz
K3QCiDO0j22v4kLOL9CurtaHY3mYY8VdI2CzGdmJmXoHJCT5D4mAtJeFJK/ENSRv
2VTZ458rB0WFTE/HCujmn8BhLbwszZhb9i+r9c+sZ5ruQ4m2D12wy2QDnxLepxkw
SqAQRRW5uOWIknOFgU2l6Xs6dvQtxIuhyr2oqpNJpcqtMpJeMZd82mEXvKJ35top
YGKaJUkIx5dUUxwPkMTw12Efo1hx4ZpAqZP3p2SSsC7Je2ZnojaW/QV3aBdjlH+k
+fh+aAVwQDYoKEbR5DVySQvAHt8Ethiccee6rpDOeBKuvhzvSZgPag2JxdOEE2Vn
T+mTVyUfo4mvHo3JA7tAVukfDoQzkUvWZS0u1QpTFnJLJbJ1ccmvMGKk7qgPUlAK
33EaDWc3tCAzZwiwNWMl/owpXSIcCxQkwjQSvRLh1Hp7HxP84WZ4W9KHkAmu3L0s
EBShJM6g7SObAgeUBJaE5yvjQSQdmc+mABP573+0VdaC1K4HhxWFnVrpFyEV2Aj0
hENGusnsOwCFqrpUgKqkcOS7YgFNDaDAGcwJHuG6KtQkH6uzX8Z/VaZfxCdDRRWk
TrwtHsHpHuBRCPI+o5Wef4TckPPG2mGwAsa1N6emruoxaekQS4yKLzHGCrECcMeR
0cjLRcsN38yqvwB470jWe1Mcol0C7+IkYwW4+F90GIqU+HaLEVtof3LYnDhk4i0q
YCFcfVAIuEvtBTOW/kOla3M2daazpsEbUpIhVtqcRh64k9KQaR9gyr+9hv9jd2mO
hu3os+YjNXy1kXepy2NKL1qcvxGARuk0slfkM+re4vN16MOPFPQynpuE/mGYutUD
8FTQmxqDRYirW+Puv5PGlBrBvRdEwMAjNHbDG6oHI3/gso5XGZ98tIQXuy+8jeTI
pL8nUiVARkDmibK8h9cbudxCrSvy7rhPinvxuoM1uAksoQSWSEue5k2usvX68tz6
3HhAyfLwAlr+i5a/r8HcSpDFLl8DHGK/oaFJvImUEIwCvDOLg5slyP4kXdx6Mb/I
GCtCB/m4ac2QNvlWcwdIgA2QfecevH9gfxoabz4KORqvFl0P8YZIhM3IC/c3W5Pd
T/uFAgnkOloxy9kB7xe9vCs36SvSmWmMgCCU/2loek55B0XD4olAt15vO1VbBTDY
BP1m0FWVnhmrWwWZBFrmJn32rpPRMPbgcz1uEhz0+gjN9z+dBWOz3vBp3lt+sspP
qbfRcXmkzwyMxWFofblKy2qVC4JaxtRgc/mGw5afCUSdjPQh7jYbpPBK9Ng42hpa
xCIZ4Uo3d/u1UexG2BKpNE9U6GQUNtjvu650rvz0xVp0wzZ4pRZTyXyORod2el48
kmS7iToa0I+P9sVqFY+GdrMWWX1/+r3pAjOG5Gff34nX5hn0L4N8FCH3HtqmAO5t
PDIdCldpUp6PCGmnfq+rk8KeP9xH2GSTJ4wIXQazf3fttDjF5wnzGjThPCdT7d+j
P+G1xmJM7Z67s+qfEEq4aWQmnvbI7ciyDX80Dug747H+UTiWZcCwfzvQSVzE7Hb3
65P1MoTh1ma3ssBxKAccHQpmxg+H3xaqqvtEO/9zB5n5guYK8aVtWGlBE1Sk9O+r
pTNe85L+4gMDQr/g796ox0o1wllw1yLnCbQqiptoY8NW2ssbQA6dYKH5LzrMT+WC
Gjr54p8Xj9hhudJ+0mxSeVL9Rp1i3dYpaKDAU6oCJQF0jOwBYXyd5v0Xt8AnaYt7
AHJHJFCT6BrEEgZt8qDPvUZScD0s46s29r7nBgPdLyKOTow3U7SMBePFqzdnvwcp
qV6GgBTeNDrzM4lU1ookXt32XaGhIowmtSA6Lm4ZARYtZIoffo/KIPHajqlaaX/r
pbl9qiXoCEg9QzWlBrOeYu2pPrQrambWEeNKGrMj9CgbEtqTke7W/M6IUZOVetYW
vIkBcP13ulGLIRLdCOFOqpqrt8yms//U2nmmFjZSRiy4sWRQW45uh7wwe7Ra+ty7
Bu/h/OzwhSrEwFbvV6pqVcmbMUxjjmkENpMAuH20L7ft8kKKM4/+i4qcq1iY3/0s
UztJVvZtPdd8TpT9P5ixmPotuqrkUx9SaVvOqRuLznHIXc+Wu4zSYHE0otBY0TJG
Ej1NTgU5A7ZNP9raO+nVkMBMuYKXaJtmtkUbf+QDV3NUBMd2pvNzyTptGmbzMJAz
0quZ1Gzb1gxQnGopMuuECV+vFhefHWNz2ZTf3+X7DbqSvvxWVqidxMfP/dn/18ht
etzdiTgIk8Q8QpOnUSK0S+dEf0EwWYg3iPbeElmdRa6nlvB8Xza2S036dLhEPeRH
KWWigA/I7CMW4awgUnIScOYByvgaJAh4p563Vx9OrRIlVnhJn2HysMGAB5faoO0d
D/ZaAXD55zFtFqwcTztmr83zYIv1f9/RYFnNIXzl0fCAdDXw53caoFtSlq0rFHhB
U3kstMWDkNbCKS9oqmYyMFVw1IrQnFn0R8fs/c+UiOmFGK7KGd0oE2XWcNUDEba7
ISzyuw5jI2CNBDf8HZQai6LFJAjKuus+m9+bJlwAX4QeoKsCy2q/7O8XAkzD3Vb+
9PaWsdI+OMdve0Oo4WfwuFYqvYJSWIe5trIb4brs7zB75wzXeEVKeRco7dGG2GqS
mOCX9G9zEZEYMCVhmdCYfYjGjET4G1yMawCnvXsQGF/QXW/YsYhccS2FirRyASBF
94pUP6T4XHTdsTYhLSYDXAU91ME5ppviNQz4baFhh5xYLGIiHHsj4F0UAnD16xfR
xM/XK67RWbqOCG1FoI/YWbrkabZZUm66A/U5uoiYXCM5IbnMzp2vKEuTfrHDZ6JH
WnKfEAuWcgGdn/NQAEMufn+fR6xPrWDRvI51FmeG1KEUcZUfIpzqKfJk2YhXwlDq
N94eJau/LtBYoXWqI7M1Bs0mYOlFeaPVS+MZFEeeRxKuhhNvzAuc/ss292KdCaOu
Lo1E4eN6lbEOdwYyvCR7mL0fKN2rceGnNMD2IzfUleYlMEnCxSCfMYUdptQVd+bP
E+PiA2qWI9lPk8tvb1BW2hv+/EU3QepBPcJ9HwfaDdgljMw4a1KCN7qzqJJvdB9n
n8vsCdbh1BjfkpUdgE9vsl/PWRmiYMgj8qxHffnvfNjMQEnGHiyIWC9hNY9Gqm9W
wgXpJHX2Dk/QBekkZpcDJwuusNRa4sw7vqeEz7FHOePkhNQd9vfOzGhQoTOG1QS6
907SZEImq+P1F0Lnrz4yPGhyodNhRQvnCNZqwLASE94YFrxztr6dNa1gCazGo699
SR/OjyMmLZ6G6zAwEqc6L/16hBo+AEZ2s1Ps2WmVIr/+ETah7KO5yh7KK1QB2kXS
JRDiVJT+m2OVp9tQ1JCZNsl0cC2GOqy9hZ7UofeIUk/OOFzmn6ZXmjL53XFpPrQ7
06hzZabltyYcyOOIOJ6URnXPlVN/Mx+hpDXkePCq3hz9Kmi7g06GnzalHqcfiTtd
8cMJvS07SfW3t+EoxJPY+8NToy/OrRJKu9tp/pOkIXckDQT5cEbVeuFfMfkOtmnM
xC4FSJSnS2r6zhATi4ZrXkohc+VIiahcM8TZ2581E8bravwwrY+Lw+PdoRDdrQJC
pRULZRowzLlqg822g0q8pGFt7rYhGBvnAto+aVqooWdbHXJr5vc0XJ+nsoJ0XNCf
1fmwFVFMvNud4T3e3x3cdUAVKtAEKwNbBPp2y0Ec4hgAYVahNNmV2DsCDPLhXe9X
MREbttww40NaoJO+DRNoZhv7/gPOPUH3xmjWs7q+aqUzSBeY9UoyaV/ukYCS5vPw
AZ7uR/8jD7PbSobOeFRqbI5R5OFESDx2HH7FKjI+w/9hiKla497jPSLWD5LMVbz7
xQzqGtCm5BMSeQ7KKnkRb3pSd8HP22IXW/k2kfXjD+yJQ9rO4+n50GAfLDTj7+TI
48JF3QGeOyBzaYGBIVJ2V4IOyZlCWdH69h8d/ZEdo0zyBjhFUE/LI3/TnGEDoNYL
rmm1YzNMeL2+5ogxSfFSBLiXLbTAKfdIJIE5nXU/ZzhreDrd0MwDHCJrzx89HWED
fcALV8SrIfAOBniJ10At52iBhVBhcD9vtO6QU92+5FQH+FYPtficvV3n5tyBadMk
2G7kdBwMJ5nmX5OBAhp668XsvqO4OSEkgwCigTOl2ECmp98LMi+7DbI7ORs8LxKn
EB4EZVGl3B8/QAdj5Ydcywl/6BbxtKJHndfQAIMLZ1xlL8WIUWNknqFyb122FLFy
1r5vmATmwbNEcgXQxeQbspFtQzbW/IEKLptswoKv+ecPZ2BmNQJnW1693/pidHS0
4Anw3ninZxSbP1jQsyLJBTTIH88pt0JKbPEaeJ/uRfA68/ErTg2Nkspn0m0neXlE
tSnN3aJjQvs9TRqwwjBxlU2hNtjMXN1n/CseHpcJi8sRIVBVXBRLlZtXx0r1M5Nv
SF6UZpjc4M/Wdh+ph9E5WJqKvyIEdEoHi9LrJ8u8UjSvOyXoYLCkpTdQNAAk+SJ8
/NO+BQJrZEz7mC2vihBSbb9T40LhRgWOdqYI5jRqVhvhg2sHp6eySVH55jkNFj5h
tjxVX9ddokBcNMacT+atQc2VWnApLdoucb/UU7/xcEpzK4VbHAlHESJJSKkMsonk
qREiG12VTd5gE3t+jiA2T37aTcqebViKC4QQvvujauF8GsxAga8zHTdaYxz2K/Jn
+qHxlRpwUJYjNQq5KiAY1vOzTUU76/dexd7BZ4Kv8aK/X4Mej4B7KdsYBn7b3B8Y
KbXZeXdxf7EHbKZvQG3Df1NllrP2jA8ajYPjfXhqQ6VPbe07kkoMO/sLIRDJpjHT
Hl2XTutr5rXmgvAsa23G0nEBF0UExEzCiSIr2By0PuOMF4aS+SKArkocU7AKJha7
Lr+DG4IePEHVRSnW3S5qfHUJZNpsQAQrCtdd7oKYIMIdGy9F5McWOasuwTyJDV8R
dkjIcdtx6kIgaruewMIDBb1BpLoZrpDSno1QxJbj4i/5tDuJZLqjIeKZRHL9SM0Z
Wr+MKR64sc3MF0mrY8NxDW0BW38zoop7Bdt7vyU1xZ4cnymi7JjdtTn7d52kz/x+
QvwQlgEMdTTy320sD5qUoK+ketrfdWadjNhSQcw8FOgD41xoK0Rvds1jb+TJuiN+
+3XuAhI1sJrJ609vPNksYppPn1lGjfwl9rUOzcCcLuEBUTcf2gsovMoo8e9a09HO
lrXlMuVnwilMxBlcdtvPMJGzPvSTMOVw0ihGIOtHwG/ytTG0K+BcnlSd5ysJRzh5
IpJh80uojw4iQIqhsYXD26apSmyIw3wl1m1ZxyqSN4Dkb2CYj5YrICUqoFlWs9dZ
VxsyC4DPMmzKDHNLXK2BrBq218SZPdBLTs3ZPOuT09dVvEsw+BuFg+SeUJYP9tQH
xD/cSj/N0qKhHO2/f+rhD71a/6EFrto5wpj0+QckuzjoNYXm14ZYUSSs0ABKKazE
a7AYwGCwiOezLW83kXtOaDyXNKKW657nEzzhZFSxwMWVujypbZhSlmZuWvo5aih7
nFIvf8eSiM5Y2KnMVktsMVRP7uU+tWZ8Tkuj0JM9bdunTcCVXtNKHjsaJb8IEXuS
tfDsRRbagcn4hmGchNjRz+LWNTi3z4T6DyJNU4o+9xgBnccRz7NflW3vXe4S+YCj
hX9vkUmj37XmESxEozBM0sK8WS0WdwmUrbq2ydVI9NXbPqGD4E3MWDuDV+THxjag
igLkcLywtztdknOIMVHI1Sy72X2vFJQK+eVEkNDI03SDrfPhIv4nU8XPQBGXm+fA
LnKDZyfqjCDKTP4/7BBNjkFezFAPpgGa8NHHZRVhbMX+juuuUZ0C3CzOiLMnRkLK
L5uwyKxZH65GQ2RMcwYQLf25k0zQVuhCAzonAMKuJpMobTAFwDBsz64Rd7FAAdZ4
5Avszu6/7xChSPo4ns58Uv4cT+AXu+2Q0BAn9cXZNUP4RZLmVwtzP7N6LOK/ylzJ
kgWMRVITjgVYUrudpUK6oiIUQiFicqG2wkRsqacyY96A+2WFR2YMMANG3+kI+c1O
5p40/+bUeq24Cs6YMYY6lCSMK0Hy5H4C0uGBBbsYNlGxrCpLHQFTO1dR2JOqpjql
1BKdWYuUgUF+w9rn9K4UgoIyQioojq1GWbUFWx5cVa5Z+Zw4pHxkAqADFAV0P6I2
AcH06Rq5B4+ks2gRKksSsXvarpX9FS0ndAWHN+oFc7A208wSeTOstFlq//JFoGDt
TpY974orPsI4JnpdYKGqqsF9sm5fJMySGF5NJBpOFSXQ2C/laf23eAiVNLtyqVCK
oPoPEP0B/BKI4uRtdYGbDcyyH5IT6IJW7adOkzuTyjOSVqvOFizZLKB4lzfywCzr
IHCX2bEdwuaPTFNpRNiwphGO3T+k8k4GnIEnOvuDHjDAJt9hIKB1R0yFrBXGucrK
Ark+rRAFCftF9bqJjMccLlWFlQgLOFOwxYkJzq82FyuO5IoDOV7PEQALj19lZWDh
vZc9wBQiqxVQqY76Nya6DHvaop4KVmtdw0nF1p83hErG93lQcxkueSrSPbq53wkf
I9E0wmpIWlyj5UQ00/llToVMLLjhCvz6FjggiK75aqrIUUG3DAIiv5WBHNU5ohB2
Nt4Q5BSA8uhBmx6iZg8EAM7i2EZT1y4FoJ2rsitx3bcNbfPh/Z9yu9d/hsraQ8Pz
spAPktSNao5HoqglELI2OnfZtdD5NV2T76ns4LV7ucQUkF+NijKZlIsibQLPgKxB
kV+SrCTeIkb8wDyPuAWS59IRW9bvfEFGpO5p+Fo/DpKnbdNhX0CZgXSP6AzxNlS2
731D3pVYRUXYul/UEvb62EpnjVXb9dmGi1Sjf6g5vBpjY0g0OpuEy4fFZDFIVjVA
09T6VM2bsym4Z9UhYx3UZ527h6jDux3rlJyRDI9dsvNNJW1up+lWGpDxefsk2dNg
nAtXjdN2FtdJu+KNmK4c06jIW/JEfdERoS5LuIYhYVquxCIlIz27AgtflEE/EF8w
WzyWexaAkp9DSH7Tq66twAiSte4qV4tqy1ZS8GvyeLzqZp5hKHjOxN7AdBooC+3L
z8+cW9GrUdj/bBc3LmTwEnvkWEUwNgg5ozpctzfQw8PHwQSEnzrO8Mkm8CMrJcgN
FnKSjhiGcCj7AKqHzhZSlvSzrF8waAQrZUgoCkOeG96ucFB7rGnMbLFS4qAZQmMa
4P2Ay82chgD/+Lnz3Z7vmn19UmTI02KorcB0hPDxldnW6BohWiWKLyjvcVZGMwi7
x4HLXEXm0coSMai4oZgLyr+94zF2xl7WZGIL6TwebAmbUF7Xd9rLq3RCjO+S2tao
MczpMr6aM2HmhCMmDd4hJ7lxOlIVQgG0/o6ubfvrA6v9olUqcRdMdlI+UZlSIhT5
z+SWBouYY2PCdBMNfV2lqtUjubYiVngGZihR8jlQgxuYLCHrksSvjbw/xNHjA/B4
UprhtsnUYPYLViISkMGlxbOf8MjZ+Zd8yq5K7AZowPKICd8jLYchLbGky8Jb62hd
51a+gL+iSypS9cKblhuy8HShWa2yWOof8YwwbLlllfhpBD56syg27URYlZyjZU54
JN6rlh7U6fN64cEtNesC5aaI3XPb68fZK0FBWfCjIP0eF5ceGq26CbzEyBafZQKN
zSVB1fgVT4rdWHFg4EvfFwr0lOUbsZNR4O5EEsn2PPG45hyK+eB0bRBaNDqsL1mG
GGcbUnkS0jP4CaE50O67C+TwLWR9Ew9oH6fOZNZ1xrxgRfEp1mYHItmBv7gRj1xL
e7ct1NCKfec6XL7oh4d9e1RMt3bpPGRJI7urP5MYJZ1iLcn9ZwalMAKOfddhYzJk
0G4k0unV0fC5L7q/qY6rFnYHJ/lVy6YZ2P7/LXoHzVbPYKN21r6E2TfqklAXT61Q
R4YQjDQMcTCjaE9GDZf5v5F96utVl4LQa266dP3JDWDazjqKnD332xBzv/9saulC
tODtvbpqFP++V7arRnHKrqtcnN5Gtqt72tFYzhDPmWgkYyeOrRX/RVCKThH2Le5m
20UUo+bMywagw/QgpPxcm35saSdjnK6XkyKCfCOBRrH21nf3oVYXQo+AS6uqDXiD
95MnUSuNKg58TE59Dd4eCvvzB0eQB8dvHjPyIoZCrCrFQAI1CRnigBo47hoRjGgD
abFoGFLBON282LFOMgD4HNeYo9Y7WtvZ4x/4YqxWhOJGkiRS8/EwVLiagZXbwsXx
UdhZemckGWabeU0fvYVIrncGo89Sk/bqHk/UdWP36WPck+/a/qShJzc3YmwZ6gLH
m816n4431qUSTop30k005hJ+8k9Lx4kxmxzGcH+8JY5jt1/PSSz3SqHn6YkJ6IUg
VVdZ9yUTzOlrQcxPXg9wYyOPBG9rIQrxC10SqlT7CyL7h1t9yZ9s3SskwPMlzWdB
7v+MeTeLNFcdXTXQbFRiO9VfOmvuRGtBf7Z9qS/Q3rH3DuCwEriM4rDSXOfIUENT
vWu3cslpc5yQZVwq6PE0zHqctjXyQd7yYv5s+f5PeZ3IBTfvC0SCWHdavCIhJKm1
Poyc31o7IHw4yQnwy62Ztj4WL9D6JevDZ2MRpoTXX3KtY3yXT4W9WK8xW+tn3SWf
ZcjcyHWMdXlOuIU7CU4xiCDPLVDSVCpTx/XJpAY3KKQ8ewn3+VwrXJi13aPM1N24
8NsRn7eWOOewdlqkzYNdRVHlxqXe6MBXgbvrUd1F2Z2lRz1IU1kbr/zMNuvp8KF7
kNlj85euBgc95MKFL8ZUiZR2C++fgu0umGgoz2iwN5J9mkYRZOftLQmc0RjdacFw
GgTz65eATSGsciB6HXo821E83W9a8MJVI3vDiUvQsyK3ZIvFfCY1UdusDcp3gQIP
1URpfkEbH/rPSJTmDdPxNNNmfKmOsDGt2Tn+AUzb2h5JdK4RBWtYkzj6h+Una6TZ
8SRxBEd/k4fQtK9uLcgsz6y7DMAvCHHNa/l1h6L0k7Z4IqWGer8vCXx/rVZehqyg
tCSZHge6Lt4UD7gqyAozp+P6RIFsnsOBBqiEA3AoDEon8o9CUfsy0Pms17JmxatX
hL3tzFaJGwI0jFy2+YhtH+dBDMSonarK7XMJ9BfA6FLFQJppaGSPyC2t7PzQ3mDO
G8eE4fjCXk049YVd5+JnghpF2Im5vOShcecd1ohnbpInDPSVlgZ9Sci/r/7uBVxn
SAr3y9/g6IMQ++nGavSfDP/b42YR3YGYkL5WfWRdmMKprGyAIyVDmotX+IDKED8n
1IUtB+eSKFLOTZZPxQjiiEZ7pRCxscFQrLopkwRTcE7hsreUHa+eWtiLMYtNFeDJ
KwsYT4lqTLkPe3HNxhUeNu6q/U0xwF8cOvp5LxkyAQL3Q8kvHZIkugbxk8B4M6tj
dzeSeHgK6cEDTi1wXfLf8fT7GK/3v0FSlQF1HQoyDz3wTgrj8M2raKjiY0SiAS/M
QFy/1fHYMNd0SutP6JvVtrkE6bJ0HiVcsj97JrRL3184cPEZhfT3c39AfSWbFxS1
BFRdbCqhIjhXU2ePD6zMwCYG1xNiyX4cRZdSgMryS8EwpjpQN1l1EGS+bSv/jMSv
1Dwc6w1nnxbR0zwFPY3rEXHjYrUqFW8+PWXmiDchqL383wNwAjVuOLmKm9tbBQvY
GCOSz5exQ3OuCAaRhxUZHLppXCc4ENgOPdz0IW9D+oj1oqmDbcDtIOWKhy2s0pga
ld7bJ28rG1DO7yQD7vhP+qxuYm0CFC476Nx1X54tp/T3bOv6MXm8jPcGaM0qnTlA
K+nGFysm9g/apHqHnk6+Fu1NEVXvMNuiYrQ8SGvx8JL09L6zyXW9AU7peo+y8Vyy
nn8JKYSeIwtb4aJYv2mhROkbheSZ4UvQbNMsd6pMY+t/TjIS43n1GHct/DTJH3aG
L0HbSqlUuIhhD0X0m9MM8XPIU5B+2iVkTIQGwJzgQGm/qve357hqM3KWHdeo67bt
ZW/jEnAvfRtr4ukC4WTaI0M6FbGyloZ+JhOoKXVlon6Rd4HfsKPFJinnADyN6qW5
UM/WLmuh49B38P9uqaTNocFlpOSmFZIrpMDLXXioatWjyC2SoujYgKg1KEp8ru+6
0gI8PyJjzL6qAoZyGq7jRER19fMN8CEMWLeEi+MkHtK807AuNwvPCvwbouc7qOhz
G8LOVZOfdtE/EXeG2O+nQXmNml/3fgjIesyy/FaE0CCQVAuKtNw3YgAOtV6pez3S
MbXfq4oD/jnEoaRijndumLwe1H2GPpvDI7z+LVthKGnw/PUQCDDEk51/gCf6Uav6
xDn1r1POCEH9r60XnQoRCWUgSNxNylWI81x/LSamPZL8pkQW0lsMGr9g4oe4MJhn
5w3w0zp4tPODKIRhVet/eFEutKVfJ1+pn8I5kC7sqDCsHp4P0kwQlFjgxZGDKPHM
SmvOQyPMwAPQiG97olaz4E3xIwwgFfLbrRlym9nEBQ/ND86sHzuhcXo0qf4rvdze
oTgtDC9LmIofFCKDgVYTb7/KDfQ02nxJOT6AKYFLfRnyaw7n3rsNMbxIZ096L5/D
93Vs6wE5a6h9PSMucVNuF3HNS8GCOK31cPZ06Dly/+KswWmx/dFK7AGCVoe/SACz
vTz4Ek4qlNWnzPXuGTGiuSATpd01UYqDZSoLc1a+uQOfaQsOg6FYqd/faPW+nSd/
6kSuztmGh3jgsr8Tp8v2WAfBP2DzTLIc3D7LrU/K5rckac5EBe238valVN92itku
AhnERbqSvhSWpAQJZpS6QWBi63Dgyf43qMVAn4rEBPoSFH6N0Sxr90WA4wGu1+Q/
kMgXbTHErRBsH1c+xXZEOo4AdCjpkeSsaCLqDZlK4XZQ8ImITrPVQZ7tYTFcACDs
UZVPUkHrQBUCu7WahOojNRJmPxJA5Hv2x6XQxQzth0cXD8GxHdN7eNRn/awfcFPN
8+XPnU0n3LZxMuG+XC48sYasq9et0t24qqnvRtZ70pQS4DQGeKa8S2vuateFj40i
TuqIVbmTURdplq1iCS9sTKRHsxAkUInUBLtERVXUuaPLPrPx+mgUZTTVK8ToGpOC
qltEXi49fwd5H992b9HqWDrH1XRhPqQJgE82Y7OWvhGPZk92f8sflTKnIiZir7xC
kkJwoN6MarbvDVRzVMHY+kxLLAOAplFxYexNei22kEj+t7xw66l+oeeWQHgqZdhB
Jiu/4a0VIJNIz1It7qCSu+9+6N4aFs7BG/dzi48THm+J6QsJheKlQOus62ksHwpc
wTJNxpbkJJk8BLw9Er1gJc9nVazUcDtDo/F6PgN24wSomHTeOk8MiK9HnaVjf50o
0yfbyIJ9/02ezVDZN/45NXb5E4JycBl4a6wjSrx8fE75YEaMAcm5jWWT+Dd74tgg
E1u2PbjVVv8ResQSGLGsu4GFbS45AwQUVvGhnj8RVE1GDFwjJlNc1E905nRPHpg8
KR74qFv5/9MflaOTunpEAKVLnrB8jzJh0wcyu6atZ/jpaMjXHrOTCv7DqqlyI93n
ebwwIG0StNmT/yWfg6W0oXwsgWMZRqIUxqxXkPwLOENId11YgHQOvZxRXIHSUL0N
CMoyKYQgf0LLJs1Uyq00JLq1MIrF42kDFFJeH6SI1+pCxVi4XlvPZFAdtNptx2Aw
lmHbEgvHu6P1Up+kqJbm3voPLhEphFlLp4lL7Iqcx3prasINTY2Cf1o7LTDyCUB4
Mto0ZfeoKtzcmUxpi93f6oYBLkY/92R9qfmRL0jqYaJ/ppsJva9OD4ycwPjdxGem
+3NcyZ81/PMsRpHYhrDn+mGiZYGkbYib8lKF7lAsD/GIuUdLf507ywbPqoktKjjM
RtKncD8PgU36+wwO7rrxieOa0FiuW8sP8dwvwgCqBVoYoKJurpLN7zsW1QzLihFp
9K/54aJfvPkqPeGk8x3NNUebfopq2Tf4eOrLHjAKMljNIIYLb0gJq54ds6jkmDTG
21voCGpbZ1feHa/pk6v8d/5WA1TyQ0F20HGG3S399Jkp3J+0Inb+79QOOEseJBkc
KpDB0XkpGZkeaTs6WnwaNpLz/seidm/yynApRRixZJ7ntqktgzQX+PtMWSpo5r9A
lmF9fCwvyIXUg84pm2bfWO7LQ8us/qh+0mPoWwL20J8NQFhHFzFnSbbCYErnyOkY
5oEH0HTxRLq1JqAvvlO8Xv2yEGAUtMNfnnsvy8mErgFm8dlESCquznRIbhht8fUz
L+79kTucX6Snyx9OoAuAQgaPg3HoAmJsgYWDjOyIR+BdWilmFEvrM2RIl/KaAAH0
kRpDZBq06AeTUty4zPbVqKhiklzVoLyS5K+1LlGEyrCNcQFs45xz8D3pKVTEccjJ
O1VtfAO1yy99ZReIcuTO3+UKyJW4V+XuXpomBdu5xLXdvBQtoQ0TKz0p79kN11uI
1GgKcsC6PsG8LzyBxH5XflGlE6HdE0CJKAfelFGOcUY7omW101d0zKIugC9cZRM/
6d56r1rDHWXBnenoN5BTZCmTBpCi6XTMcnfckvy8sXw4Lya8CPsSmwSxRLmSc0PD
BsZKpS5S8YuyfkxzNueVgGRrD7SN3frXmVIEVtrQkq+6rev3Xse44JkTmFjjtrG9
7TAoK/C5IH9qmth7pkc8rYg2Vu0hb+3rU1xRKmKAZn4ZowcnFQgqOq8VKU2egYt7
K7DgaA6VPV2bolRi+laYm6skDyYaBg5ocbRNHrjchw/oPJXhctYiiWn8JNXKcL/P
MjeA0LYk0uhWxpQyu/0n4tpxr5Fzpoz85YDNTYoZAiX8MifbLM+4RxSOUSLmktzV
NmshLh1Dk2Xl9ukQvV5c2+arty2G7cG0juADzr/GNZS4eTXmCzaE8voG0BRNywji
2nWJpNQhQCC4VEpozmBvu+LKUoKokzTlEPdqL0sJNjq2e+Jm3ek+OwYpVTVccYub
HxEOnIiyiUkHArQflJhNT8CMqc1F4bX2jTzoKTf5PS4Ll8vY3uPRTQVD71lLsqXS
jblhDbtWSEzl1ZO6mYV6TCr0d5bScOq5k8TFdsEXbIlK3TFsZzLvkpcwul1nApoE
Me0obTMuiAxkWIf1LhxuIzgflTTzpqgGOqH1rs8VU0ce101E1Uo0/2s7O60j2uGh
rnzp2T1kuUT7/E/3gi7ftL3Rm6A0sunNEhT6WJW/eLAQqAqrFzzNNULL2Ve+MALV
odE3o/erwxWrLgNZXNlwWUaYQWTBUt1ZkROkPHayrZ6na1uN7y5O7oxUcvAMeWz3
dqviB0sXpmXdM4OhDXLRHXz/lCbQ9lNhoKxXi16J4v/mRhVbc05+ZwHtMRkftJ8v
pmAVUMX6l451GuyZAcTfjCSOhE14qRwghXbcZV+FFJ9R4NH0sqlvMglc5Z5tH71h
xQNGdNHoVHc+lskGAWJvLhFG2gHZDnFheCU9CQ9dO8yj05/UHgbFXpVjusMHKx8P
mAO2ypKb0A64tnVFA6cU+8MwyjnABLLce2rQddFL/Mj854hAA3wl2IAfptmDkdgr
PwXDbX7uDf4QSz/+7/SdU3TDLKqZS3rM9PSQgYq4ICjvhY1zJruRb4EjWLdzC01g
0U/L+vwEM62mhbGvBxn+nQr+0E7cRQfVumCV6K72mOueTGYMLTBXMU07uNJ9sBUS
LSx8KQpfLsWOcr63K2ZE0s9EaFFh42RNS7WAOx8pao1D2qCG5iqrqPVKGYqYgC17
5gmiuXx845Y0AhkqUjBFZQg6csexGvqJYbIppPZHO8R+k8rsZrNhvUV2UBb/LrjJ
hUe7kYV45GpNYlYgoJS4Bc4Y+smK1n2i+8fXTQ40AXA2nE30YLniGTx2hMqO/o0K
zZfj8TizvSD0tBeO62tcMEVeTLgnBY4xC/kiDC/DJhhasnPnx09j5d6Uh6oD3c79
nyBUGhKWXOEKvueQdREXcJtYMXpjruMBBAtFc7G/fNS4DrAVugBfkETySawER2Cv
c0lVsl7hpmrVWx1PfKsY5r8pkEP8x3NNp+UxQWBOUj+OdadjSSQinstVkFgGwKzT
js1krNBeUOx/chUxc6BahaNDDtysD5W5npKmfaGsnovXoGgn70fGXgrAYb21JA7Q
JbTAKXPMPN6w0htVCtd+Dj8G+qfjsF7nj2nlLYXYT+0RkOftdRve9IjulYhq736v
OGmlTAYRQx32O/JP4D9WooKiSQ8t0wFTf947tIv3FJv8LS+cvxB/ZRtG1tLD7x0L
upppnPz46C1bH8x/MT6r4Z15wGhumC/+mNhjLO1fQRGD9R39YN9CKw7DgQruRxAq
4Efbt0d5mSvOEZT6UhxEpgFBR/2IrXIyLtNE3FUkm/tu/MFmq7eA5KTc7NrgaP2L
i5eAOK4tGNizypqg8bEE6MDLJyg9kLCEJxZWGR9qiHafeuHx57/rPMAebfBBcy2j
GJs30bKm98dQpm3D8iNO6Be9qWKbAEU+RpXlTDuQyXlFtg3ilFOw0P8pWlQ0QuNB
KdQZKOaRZ4YnTvu0bFDrCd83Q4lNox+dTVk0d7moGHE8qBvU1zOalUDWPrsiOM6y
9jSN4QwOwlJ4g0TyagPC1Qlg2nzVAgIkpkI2vxS9y5hem5lInBopb2QYjZwP1Avv
/W9BOKP60wrMkXIsKQIK+Xa2mBik7Kdrrhg93PWeqM1N9HGJ2xB//SwWlsPGpURi
FkpQxSBJ7Kjl3OZAYJrw+E1hhL0ISl90KED0UiiqEbTs8LGZfWO24m52HK+9F+Dw
1eaz8pum9gJ4THVgfDLDdx6XabsVRZAosw/NINNCKb624qZXDg8T6FNbVv7UWJdv
ysm695SlkqpSLFmXvDGhPTKc4deEHlH2NUulJenZ0PZCeoCWMimCWXuboFpNQ3wx
FsVlWUI3Yc8Ls8SIRfrpYTkwrIWeT0E/XBOc3NcqxCXSxPL+YPiQWdEzkMNet1WY
DScsRiVxJoIhPiFSo1ZjJQS/W5rAkub/tbGlimMZ+T7KtpY6ms6hVPG+WZdAA69X
FZTxadY42J9P70k3qCdsuFiJ5eB+kaa/vloi8QLzUD2O07fu3PTeOcz+JpGB+pCm
nh0w0VMsSg3lGsldKiZ2b23oihf47XkZ/WmriZE6uC7Hyv8sxAkuZtBQE8UevNov
WKVIoOYQvltcZjS3a455bn6I0AtGCk5Na+49if7MpldWheyyRS1UNDB15ZhFhpdK
s92RrfXeZCQhvM4b/qp86ogaZ3CH4sYEmbWZd7nXUkkSxnUU7DXNN4USXhg+Rixj
3Q+aC17VSA+vNUsm0WTIj+iil85Qeg28qd6ZujZ3FAmS4TfTT9dV9pZLozrhVKTi
zcdBJkUvsR3vhicxxsYQPz0G3OhtSYzIoYE6Ktz0jransGSfP8+UX4J71N+46UAM
g0hSyq90oNQiC7yHrbeu01nSSfyODloQJelMiAq/Az6lbekn+tuoy2G+fV1Fcy7M
so79jfJ2Dhnih5ptQ6hLnf6iW3Drd/awiiD4c1KEmjNz/egXFhu5R5svBjpaB25L
8aHpAZ4H63uEPgQ6W8V4Jz6x4CouQtnmMDOvyjHfC0BE8N6Xd/wupnkdNWaRWYoo
gp875u9iKPgDgAPdAxJ8QihXfauCE6Qo4eLq3Z8lUj2n/VN3/4ABUdKc1bZFpoAx
+rw580tn22LUNNaLRLD8COE2b4wfrjsWpwMfSmcTC6EZjrTCaF3kqkSJ1HCaAa/3
g//K30pfvwRcXQFr27K5UWTesXMmZJZVWt/JdI04AsGGHkS2cRGvDgostncsj9g0
BsmwYvgHT5MkdZJ7B+180OlzWtPbOy9BgOrGX2XFMsGqT6HpVoFxk97u50nEOqEE
jGS1nmY6bqBkbw72USb17tj1uxKSTxmJJYZRiJj3/UfYVWkbA/WsSXlKM/turteZ
WKLqlMX/Aex7J+BNqQ91Ra3dx+iktGD65KSqj4euG1nq5BFgUdyP66Xzs2j4rpM3
V1/Ak8HlgNyj26xrriA2t+I3msAul1eaAVaewkIQqm68EstaDdf130h40vxf0dES
qP57YRuwL5kdUvtwAlUwGVBiDtsRucsRaEMuQ6IEdPpWwMARFxLFk718sINM4txn
kqAcon+ROhU1OsVRJ2mUx+zNqhS14756CFR2/4WpaEej5otqGccBrS3cv8EYkcON
IicFwsetqgR0kUoUKStpRgvCKK1yAVhv5vuI9Op12tRFcfvhTEKcD+8FF0kjN/rm
KpF4//FbpYRwH9eWKk0mRg35+cHkVS1F1sHIUwbPcyh6pFKW2uoMOnYPo8OOyFwb
5Y/1JdioAekpsK0dj67qaZGZM4U1YPUYpgz56UYqr8LBMlW8YEIGT3sJmzPOcd1G
op4dGD/zjFo2jK6QUQrgIg7RW3UMKC0XQOf1QspNeANOdskZQrsjzI68kQszsgze
dKC+Mt6Wr5NWN+2uI/BRIZfTQdtftoPS3krxpFJYWaKu7UQiLVXUGKxMxreEXOUc
ZXFcrSsg9TLybhFyV2IVpLGZOCJlu6GmGuF7BYW4tG3GS0utwqZ0wid/O0dx0ET5
MnmzVXH4sYA+93GpQzrjnZ3XSz9RIqEqJU2NkZh3lOWbjcFIemGK3yK9PB2wbxIA
+ne8TdghGY8AxAv/X1/9R6gvSIam0Bnt3zSjiGk3sbG/+437fC8r6rupUR3wCzAE
I32eLn5Fc51wXU2V4d+T1qeryS72PA5Kyd98ca7y/mESiOUC7WQr4K8i1gwZBx5z
LuBpVcAikQF5TFFFGzJYVcNFWRPmhs0vTW4AWEDaPHK03qGNjaIYFex7fPvhTORt
54IYfz3ra4zTkelaxlbgT60pcq07CC39fB4ycXQqFH/u4AWHGpwxEGF+vPrhF1eE
lQx64IKrT3z/20OKQJ6lhwssowUN3rheX88nvj5OkFFQvP2XLSQznPFnR8csAlG5
JMuoxCaNj/tUfwT+TQc/Zy4Skv4O5SXZylV1m8jLGqSRpk+ilkiolil2psmlB5ai
Jrp3/Gy0tdFu+MNMt2uppp0FaAriDKbWRIQUUjFZhKw1rqzKN5IOAOxQGNkenB4P
gtmLyCMoubRRRyhfzNrG0i7okx6Qol2z83OtXIhmVpYOzoPXZe+VpS7sA66EdUpU
bKYXwkJxAsHxUDqID2W84xmTatlrhOQnE2tdx9zjwT5mcAq2tLD1H5QbnTgKJLfR
ExHVrAXAvMFfwOD1CPhc9spanMCbmVB3fbAswSQ019e1SC8p/d94j5HgDFmqYSzM
CzAIPCz4e4IqOb7zLY4O/VwhX+4G4Mr1qijhnD4KX0rtbQyRQ/GwXn/84i2Uidgw
fvB4KBn+nvB0z8wniBRUJ2OPoU6sZGAKhFvYiZJu4slxfUj+vKRm+oLLkR0zhr6U
CYKw4CS4YXFFSDV+Afk5waFH0aD4Jr5hLU5JT2FgGdcYsJ9bsKiyOmjZBH9EDqgr
2n5ws8dULhaTLtuGU1rbR2a80O2Ld7JgdM7xloC6SLbkNIy8z20OKBUnqdL0mpOs
W6+eKODJ2EjjDbcBakR+zvhUtSB4cIeibKRL49yICbO8LhB4hCmpnruZZ+ZiDBMd
ucKbaCIHnSIn3mHsSAt78Sfz9WtjrMoMxUQcEfZBF5pLvk1TpFCs6gRvJ5VvgVxm
xRCwGnrrNt4Dx7jp6YHSqOb5gzh4Fcx87K6TRYNjv3zWzxNPif75eROmBOfcMufB
m/LCs+Z72PGBDav/guZzYnjM9tWxwlMUFcgrGo8iO2ZJBAARX/8vpzYpzAHjJKri
igGe7T9RuPtQ+MpJcGJuwLb5ecbys2t0lvNK0lbmsbx5JrFNy3bRTpQv7RjVe2eM
vSe0EhNFRygCm01CID1D7Y82FYCyUFo/mMNF5/o2nUwtReeh5teSdU5TfjNUZ0gw
o5XM4l6WZp2gfPhoVbFecvk73vgQJ8GSla1V1t+0O4YJpe/qF+bp2A1YPnYi8/wv
/lfl1ge3EL+cnEWKdFinSb2eT/6ld0kLkKMDT8EhwQUNaBBRMZrP4aOh0RxqP+GA
BRqVY472RiB9gQCU1wKoeUkB5aWwsZgKNLhJUW21tC78K5Yd6WeKIsLPnHwJO98V
aMgo9iGCpQWFpwCf584FTtwoZ3FBYsmt8nNR1WbvRL8xogkAO6kVY3LBC4NT9UTj
W7LL6c/h5nKJUYOoz7/zSbNH3IF3z3LJgpFPGjttvWo/MxYrhogeOt8oeHDzgKNG
lIMZm5eyc1ahE4UaidE/jAkEPzYcRcOaoLEb74M/gviE+bu7VtoBo4qE9vK2Vsx/
NqSJSVcD/fnNT8X2BL9o8jrCVrEp3SoIZB591adXadgwhBIpu/N8bg+YRVu1xIxp
xKS+jMFZV0QW3krfOHfYX08AEeC7MnegHTqoz+DqarMC/RZZWOcAdJqTUuBu3oGO
dOvL0G+qvuCUoUBH8C4Fz2Pf6kAbmS1iNUkmgULd9e50J5EckIPcgVmbVGZtWrEE
+KNScfnBYbxF4Z6QD27hhrCVjfqjGN3QmNzr7k0U0WycQyq2V5heIttVjMHTuYoS
fI5rgSAKGk15LbmDiXZ3TJq9794qBvREv/d5t5Y4d78wjjhp6lAEYEI7dgXeHiNw
3to9n07CGkcGvtJ0qpnvtXLuM2Nbrq2RWhb14bgksQIpkj9tS08Q58nCZo9B9kyN
48HBWjouNoW//TTF+Ld8b3LRiRwFQAq4kXEDJp8HXrVk3O64PKz/ejLSAreOjwO1
R9D2wDJ4VTEXWKmu0IblcBtGa+T4/AA2blGh83JkT2INMza1u/pGByXi/N9O/OQp
vnUR1MdLiMr6RPeubTJCjOw/CZi1CvKUYwjsXwEBXqEjQqhYuG2jinBX2ezgNw+n
/wGgw1GEPszoN/A6ngVRmJnxuiOZzUNq1dPP+6w81VxU9xk2v/SFmyNPNWGN+NCy
72Qy27p4150z2EJVKGPWyxhSfqQgdFCWUAkfAVR26ybBhhrNxkRaQP9L6ZF0WRPG
DiD5wJvCz2LpETusadstnf4dq8ey54jObp5eZIxdntG7oABCV6nKkLUj/FYheopu
qOq3BnEoz7CwJGSkQUXYT8v4H5oWz1eTbLNrGanxThJEojC1YKIO4vIf0mp2kaaw
na4STDxACsM1ehsGlvr1VXc9dM5E0u3kQH4qIlf2fIurUcAcp95xbx3tvtU7QmRO
3e7fuqiVD5Th6ZuCx0ODiNiDU6ewWd3U4p2kAzL+8Gl3ombD998LhSueuxgT+MME
zZyKGF5CeSvqWTB3FjjztaLfRJpQ6yumEWrFKplap7RZBznMOtqb9PkP5TLsoXTo
37hiaVl1RZ4UrICz0a/OXCiGGGgpirYpUKiNqm2BTeeRvIazhpA8x6bOA2VqnxOw
MBSyutmQxuXD8/FtN1gnFCd+KZ7ePDI/QGmLCgQyiMIe/3LA+TsgqlOlzqW5vPjW
o0+rDCRYlNi0VJuW8jfbhic00bbrHEtSKPVFPCesU3DYLMtY1tp6flIVIo5sx5bZ
YhDFfTGRQvYZD2+im6Mhvz+cc8roAReUVcFjRE8/K7dxLB124gLTefl6aiD+o0De
CsHIt0nUb1ke7JK9eBZj8cxIkroMt5u8tMdPw1dDfRNzYFPPOEj5R11AkKWr0MPI
j/QI9xR9c/b8RDMtZ+eIfm9A63+F8fZtFhbKd9cxurI1aeijKLmuAGNq+2tRTvIV
cIu9nTImIuOqzAfkfJ9GIMYoMynWpL/xmMN3TZWWtggaRxGfkRjABgCYJxRVgLgw
mKX52ebuutZd5ZmzLC8kQIBEqnipIaPG6tffegpO2nLKUl0yhvTRTOYkutV3LYlK
bhnRObgA0RAZFr/xBzxSw5y+1qohoAN/jGAHlTAdtjoGa1irmLTqAxUleyocnpei
rAGaCoH9VItoZuzk5djwXMtZhKQNgF3XVqQ2lgUrF8SLAdE0thbZi2p8zbK+xz+o
O/dDa8pWZRuyW4xy3M0D6JrLdaioYUYyPaFqZqTIb5S/aX1b/R2IoWc9DOsbMKn0
lyY27YX2Frj8OH/PrplvJ6mvg9nIO21NYDFntm5f42E5qn7hmHTSHWgDAJXBTMAf
dOf2A6iyCMExhYSQW5iLYV93BOzozW6F6R9qaVmqMvJhJhGDCMjPvm6UAZtFiAUo
Wmx/MQyeTPSb0ObjfowosVbywvX+tdEq5MSPCa/QDkIKHZap/DGqmkKbaP1xGSwp
vEnHSjURSe0moHM+uEFis2dkTzs/demAbAGyEgiXRKgV8EX7ZOsSHfBUwLuMaJTB
w3+3ZgtPYx+lV/QXNJSgmt//IrI+AXBd/QlZUagcgwh27cXtLmsXoqhfjkMVSYOr
Ui9a+h+a/jVRMcD2fZZ4TmYTEzS5u7OvinRYcVrUtUfWPmij2cMFWVg0ISeYnsWS
DRHpsxFfmQdK8/dLEHBPlEAQso99LxvDLyB5Zuxbsk3Abq8qfve0+CrlL5xV8MK0
yNTkSKPyPNxlEiFSwm7PjkkrgMXoRDeONftP4j5AmJDZbU4J2M8eEl5uRpFHMb6p
6uSh7vo1RJMfnlisWWJ3xs/etMiOqWMTXC5e3Mb9rHwJ5NnLGMK9vn7JBaIzmja6
7ij3rVL47j/nX3xGuHYnnJwAgFjghjSCtBp2IdzzhFY5nDzkiIyoYa4Q39PDURyZ
KJd7xVDA1qffs9Q4HhPS2ThN6W9LdtF2Xd1UGGjmItJAY/DBYhqAEkqFcNvjHtP0
51XKoQdoeDrDStVxs4GG/hfWxv19d1TI3bq8ohQT1OnXmoVNRarn4Siif3bfJZMU
4vvT66VO8Ach/wstMU91Mit4maDIMdoup3OtVR4SU5MnURyRUuVX7fPTrAEcfTYM
0czGTIQ12t0pZ7R2a0Z/veu+ZentG/xDfel5I47/4g3YiJhwrKJMQRiI6hDvI/ap
wMU81CS3aX7juS1PUoA1qwBcFnlMXHk67QYB5qChd6mNqROe/4C6NryoTP1mHfNG
qmYl0Koc5TAql5bP2LSCl+o1Av8Phik7NGqXZWskpBoifOBlyqekpzxxBUwygn5J
xWg9a1V5MI92RF4EqszDSHUl/N5J+HER5tp4HX8NZTuiiZTke4hOU8F40oPSUyH6
UYHW4zqRbpqXpkH9ynDLKAgu4zF9csnWAfxqz4fD2qCR5E/qigR2lVCRizoy5QHQ
N1lzvxOmGJEUs5vB0EOl58tPLVaLZtktoKX77eOUP2WQcEp2dVbOsE1+pECe86Xv
Il3mLgIcuYFtOm7UlHRmvMcOEpIOG3N2zS8KWE2PHK82A3P+68eP9rKaOTOnGifC
Z/L97qDJGTHDyTggpRmCf/3M8bckpD33AK3D19wVAJkXtnvdxqZ3y79mWc6sVGOZ
LhLFFuyvaGTcrLUlbCV5x7mNhtvLcBG7PqwR5hKOG+z/HkcIa1TbanUljoXI/ryp
xTQC7mYyit7RAvbmj+r1VU1vK13haSpNSVvAIkusCchGmMIGpHEwjmY0si5Dy8os
BEzDiZYN4k5VwDzn9OgTDIHFeX3zFMHf+EDtkD47pf71vFsYPWZVI1udhGIB2jaD
3BbSwdLuMhZeBiSYDrtvVbExit73TUq3aEIGaZL2Tw2YcmjitjuPFtckoadtEQxh
uzo/6tk+ju5tcyEFgXApUpF2IXdBZ6pgJCLnzwQItNNb84Hd0+yQ2bGTyefWVlth
GeMPkcrSMzCvw8tQmsU+IO85WT96uzBlsmADDuYwsO7lZwHZFVgUYTzuHxMRO7Jx
3bLqEVcyG/ri8/82CPz0cumgOmpEYHWFcx5KEEUPqxN/8g86AUrDwVJdjydUfZIK
mhe9xoJLyRMRIHwuR1NAHwArI2MGl+CCWJXNI9sGLI7Ai3Nc7WMq0+XsgdKBckNS
v95OZpXbafZ1kUR2fl04ZPQ3XeEdn3l/BZreZZon4XhSXaV6M5rPzMaQ4TOMp7g5
efwzIeL6T6oby9zivpxWIMoegBssbD2walQwfEICzpOpYSWn4xZl97GmR/K/sPC5
o8uST5zwIExVtb3hwDekK9O77q2M1r9gLNQb+hBgpfYLDPcZA5EM/CqpADoVwnHs
qIbZuLEVV2eUMcGSo6T9g84esYLfgdZwZVgkiSu7tvWWWnbqoB1fIbHTKXtzYWab
rnmamZt+0tyUr+9p9svxAXBukuiTCbl97Agyc6MI4TU/i9JefsTnan/S+5sFbjLs
BnWzSPyZWRoxHXeh8AP8om7ITXviS0a8HgHbwWyDUNbk/SIiRv2W0ZlTzXXwCTse
ol94Mc1D+2p4m2dY4TIHJsyR96g4yQ3K3FZvach0l2YowIwY5BQd3jdyyMnxhJqM
bNVNY3EQWPSyQUGnyoms0O9/a1b4s0ar5w4pXefN8E1PNQaXzRK7Phz7/zUgfO6K
ZdcR9t4yGIf9k+DgvPsJr6K67qc1+ESMY9GrkW5dARJAsXHs7TBk/FwDN1D69xSs
wsqkUBde8GoePpi9fVH+4CUdtVQP+TLF1U7+mvnmK5NRlvwCTk4uvUquFpLR/OfX
rgOckz6nigHR0CwaT2CdPKp+CyWYMO29tLu1jZEKGIe1eWVwf6xv+ap4TC5nJVxG
6pHKYrUyGRyDu4INo8MBrQC4crNe3l6k/0cI23dj5tXFkse8ej0qwsr9B234ubw+
DNfyqxDwZ1NEwpP8RIoMqsdc/xfMRxVXSqpMF0t/R5PEHOXaGhhwPPQ86usC837y
uqhIwA7Ll6GtvSih9ZNERbhMiVE/H6Fh9lydqrs7N/+FVcp0pmaJX3IR+E5rJOcU
7Q3PFq1J8YCesK71j/n/sWq0Se3r9ClpUtYyGwmr/dt0MyaYEVN8HlaH3zEcgxZt
KGTxJQMQjmKxumu0b3kte05kG/VC/wYVGlezLhRffEFcDQX/L8FtSlXOxNoE+Mtn
RXzkzCSEROxFbG3vGDzdGoN3KQrAO8kaiWZgHEFy2hkTqbgo0uy2apsAh41XpovN
nV5PvpayMoVZyOnnBppjt2jMRjVcKL5fpkzPlQlgJZ4wLEiRbdtf1cCoMF+pyK2m
LjEAgAA8J7rdNKy1/IBY32jq3zuQLmpjtr/lZ+nfSFtxIWcdRR2moH/G1xwLH1Kh
OG4dcukTS/KqHCPY1LtmhuyH+Xod5WMHr5XQJqgvz4lWiGfxS3/9d7c9MRZ6TdfE
JZM9x+mVGpU89O4Ur56jcamnA/I9dJ6E1wAtUCmaj08ovx0pLWHqRlrk+NJ70AtO
Ex6c5JE1Sdmc1mEdcrOCLv6O6/M6yTf6OF5g7U7jkPdlameE5V5fC1zp1soP0kOA
yxyDcEyWCrCpPHU8WhWCovQJjTz9udeHCG/9oY+C0sf65I707fKAkHe7SXvmG1k9
3N9LlWhlKpoeR3TZ+BNBhk1rx9jpFoYPaPJkoEfk4wKW2oSzLv3dG1Cx2Fj/wVFQ
xstt8OC3MrMwJrmDVP+YeD5CZFDXgMMJ5TWnUS5eHZI/ttzB5dFvor5m5Z2UJjQn
vUzKxc6a1sdujSJYPZt3ZR2r9tz7v5THWXKHVtvosnzEL76OEpfmdJbW96V3rCIx
JrAySYRCmOYe+S1c1GZ6BTudAzu0hV12pp+jpl52w2siI9KfHfSiAnG9sZyy5DPz
0V7uEB+Fdp5KeUCxJFZu/DbFiOrBAjB3gutFp1A1rDgtzBMXW6N3P7UpTXoj+/Qq
B12fhR6JdZKheHEPCeTMAKfGh/0NNGENN9u4t/XIXonN4TdlW4oaYMLPmlrM19lO
InBs1h60gZNEQl1qwT1erJnJscsHeFdaRr/XLWTYZY+5BDdOoI8ZGUSx89RLgAsK
3PX+/WW9ni6u2WutOH6VCUV851LJVG69Fzv81LSE9UF0TL8KRNu4PWkurNd9eHf4
i3HZdpvhTqgI7o/AMsbJnaHzRtMLioYk8fVyws/KgqCHL2yuxQihSvFJaTphyZu2
tUPGATitzycWhwShdHqjUOTfMKIB/dRqPgEQTbQ8MJ6CYm5U8zAKaRQbWnmZrdIH
sNCtpzXYgyMYXPksfZbgRBWyeCshmTOQEBa/uw3Pa2wTzaL7zVY8aanegYR3mNEW
wgj8IQmlbXgInll826jHqQAcY7wk97UeZg4G3iBzyqVly1DyVT0q8gs+lb5gSLQ9
+1HMv1fWu/0re3e5p/se1dFeyOUXzoankDXZlYiK4HZLKBrJ2xR4/JeYyjB1ueub
4Y240ufT8Q9Te/BsxPGDgdlAjQvQytaA4/P8CywtDw+gF3iGqSqX7YNYmfERTZQJ
MzfHeZ5iIyJU/+0asL3VREpLe3yTyJHiHLKHKtY3ItGyKhGt8r1Lcf3/okngxa9f
hIJM3rjwSgnsw+gzjtfYUmbXUWdYqDGsSeU3aTyCrRA/Mr8PIf1/WlfyRdLTzzRX
t513k/a1kVfZWLjXnkUZGBuSfpQ4Zk6TTZGQMxSUdsaTG1vtmaGPVgo648xNIa6o
mj+1ch26YJJaWl2JHpt0cDSuwiOoru3OjHfy88PO4yOj/Ok+JOdoHU4/wCc1TGPK
q2p0r/u9hHBTQMugwCKoKL15eSS+ivGMVnII/4dUTHqQEabWzAa8PgXWxIWhnd+n
F3fUQDcg2d0ZGwGuCazaM7YaEx8mIRCyWdCD7LIqc8xqZ3PN/CYGp/moyhS21S2/
+RZahuBrcvNoe42atnD+iLRoCkD+iDXXrd2wZdVFisYLqBX/JbDR8fx3MCX1iFf3
mDuVwqO70At4m4JatP9Mxj5++DosSNmiUeulZUK7dFrKXUHqPhU1UlEUa53IdyNt
XFMCKRxcLTLZxUQtVpufO9I9fsULfs+Z+DppbI231GjIGQT3wE0QVuHGCanuMzAY
0PwEp47YWx3HW/UsoAz4cA8gOicombxWbU6wBTgLYK7Dug6b8L62IybvPbMg/Lgd
HiYsWkQjGXIL/pVRj7Jx/Ipo6DzR32o/0/6pczl565cfsHV+eVvVAx6PSLY4FMQ+
KRxhWQi5rlK71xPjldNrBdf5HiLDu3ZswCxYh9VUeVmBT9DpSq815hIYwFAxZqnC
uJh/nndphbCRGZasCZkp97KttXAfjUXSqjTbUaLW89Jeo6m3HreRejRDTgABywcS
3cnJq8hFaNzNcA99BBzhIcqHbWZ153o9NzJ6nhaOeSGm1TVEvTGnI2gkD1Sof9qm
lA0c+qyWaQDj/F1wisz0H+1b0LWdGm2AKg39DAialPF3IQds2wCyna+shQznHhE2
/WGfnfWBZNZJ8iq27pxAZLLDpZhJ/cRUR0aaa7cUfU7CbXFquJ5uXT3XLzB1YWiI
FcxNmScWjN2FcGQN239261U/6LifoRYM06gipR+lZOQ4VyUEOMVWDNSZt/ojt0yX
l4fBcKdF1cP0HT6+Ty2MygF0cLbdZhW9bTzu4o8ZKJvbFTKFaxsvm1uvKlHOYhkU
gexDljVLoC6Y4I7llcYWWyyVSay8BfO7W/Tz2E8bRkq2a0dqdTRtA7MD6YdkbgNA
LHh4oktcmzt/IpilZ8YQFW8EA9KGcaCv++x4SWMeSNJIRo2NiD9KXpsCOyVDU7h3
ISXYpuV7/n6lDyfYtx1WNazKwRugxPXY4H622yIcqjvDufNZcG/6LxagPW44QASc
eu8YTGrx37VgFt07ttotBFuKRxRO8aqfdxfyQIaq0agEjK9avmURZyvrXwjhM166
y/rmCCU75jU5npJj9xpZvFvm33dvs/4zTaKzpDBmfNOyYT26+tc8/bOzk50K4NFH
qIL4528XdsjGL8MsX+GfzZ96kYg7Xp8M4pPVV80FwVUILJ+YDNIeeErPcc/GES7B
NvMJa3jO4jdQgsZcTNt/HGnQ0QxyD8a/QbIV1wAJi1BQv92S0BlFJb8chCOyy9b8
x1nyRjaQXRqeL63+Ssd7o8HseCEQr52wuvFzEqwmgCW933zncrvwKbR1d1DqvJOt
GtHM2zyIFzBU5fE8igc29itnDdHUUV4FJe1e2sI1Yc1O1Stk29G1mN5PJUIipgUu
20yfaIdeUVd9a/4xxdr3FlhfkMtOfwJWuoqfSHEoo5BOgK3kdJuhYjQoh/2ApYYN
wbD7uXnoZuIVJhOcPvo4cDF+IHyIMCQxCEHWqDCiJh6Q7RFQnpsTIC2lc1vnrpzd
d/1vNs22Gwko4ia+49a9gZYYAHcJSTdynVxd9rawmEN+rY0nL64uT3E236dRSstE
OFcZrotpnmfNUMqOCPEMULtxNpMkKikN+aJ/ZqtAMCf+KHxrv7BnptlDXotItz77
6xa5kKejrInQ5bIFxEUCMX8t3gb6vf6f+uFIWk3wvOOOens3VjDANp5E/s/zwl0z
owFlNoxiSaL4SaYLQ4gUdtLR1R8DWiG7w36xHRxsXU+eNaJLUjI8pYNlG7vu2C/4
BmfcUMQ4O8VK8MfkG8hqWiTILg/SC5Zv7gon4Dqf7KqeYwr5ayk7znqdCykcGdW6
y5VZhcEU29e33cQLxeNDkVa61Wo2qLZHLrX02lBw8nFN4mlafep0aaMNrvWCzypB
ro5KjOkhqPRLmkiWeyB1jMrKUUzOKYDIAfTTIcSO83NNfh2Qb/saec5X7qel3mxO
IZZGcryQ8B/DimmdfTGfHCeXngEimv3K+TzGetZfZ+bf5Qqv/R1NT9FmxhAC3Dk8
40/MjO/TIVpF/fDTvnheeCSzdSgPUim+u9B5WEpYGl/SHRADPEfrqkMIf3p2TcBg
X6IR9NAh5bSwT1WvWMllWTWO6XgHPCjT3d95ywqX3tdCBybeABifzLvnyGxE7Bwp
FbuhFAQk3Cbny1yf+JKrmJojFSWjRQXD0ttc+G5d3MoNwYHUkYvN+SY+i+ftwSJZ
dUVflLuKkoxcf3l+qUI11aTUz3YybBd2nUAQb24LP1394xSEe4UAV0QhdWINwozs
3qr1ud2CpfhwlXNKAWt8Ea+gZGcrPdwVTDd0BCeAaAi4mAYHJ3pONn8hbZHOi+Yp
dkJMI5jhiL7K46WY3yz57vgXAEui3hM5Qx6MzvdYi8KJhrCKu2UTE2mOVJCAhIcn
3UBQqQz/VOyK9lm70Uc3SmhhGL01O+rmg2slGXA/TWqJsL29x99jzUDSHqfIMUvb
wmwYVxrtdgtszBTCAVX8kYVUCWgGi5PiCLRzhC1YvsUNU5tnj/gHHAMlSHxleqz8
xecgptlqreM0U3n1dkcNuMCVrhwH4O/jECdyFHtkQJzaPo/R7oEDTyqdfiRXUpxd
v4xmEiua+3vSiYAHKQ4vBbzCcNcd4Ash8T4ddLnXsaE2P+ZBI1WtXqRKd/jbIRVd
NcNLY8YlZgqpNxPl7pABazQcUStmfhz7Ex3gcHeDf7858yws9jY684SWcP6JzIVM
DcmWp2wbzRccs/bCdnzjlqtvcdwGqSO3Cn42TnysOpdY9TsT+NiUyiXa8f4sLaqg
upuZnsBX8hl1WiNfK2N3mEWtF4BynYucQpugcqdH5cH7lgnPjhLoYTeV5brfvqpe
oCEq0SizJbI/jq/aRmnSbeG06xJ/PHCaR9JHIGIlciz6DnppkLYOLB+oLrN7YzVH
UJcUb7qOVVf8GWLqhUffaQZLnu6jKZWm3Jl2HFvRKF4H//xYn8UUcHQe0UBq4/PT
Jt0bkEJ/iU07t2Dxzq/pSFIEhZ6ny/NKddIqXy7yShKaO+mbw+b8cI/ECLfCsVc8
40VXV6YaECA1/3frAZlYDzLqmrLNs420cPiZmV/7l7wgiPO3ju4lhsr8vkXZOPYQ
0PdqqyHw3zS1O46Edd006wZ51UrNUc8OoKW4KD6Qki102h6vA3fefvBOwgPz1ZrC
snLfRJN8ao9YGzRijsHlt/qY7XfMAbGDYxMq+XvEtc/0DRBZH+O22iuoyArV02om
Vo4LTvEpk45dS4g6QuFHsamUktWNz0A56rXTkoQhR32OV2kXevdR66dt/y2ZV2Q4
yu/vw00Hq6tNh/b/1LBbs/o+c3iNpf41ku911lBMtDr1KccWpPACBNR0suBiSVSu
q4tratOmnaueGiYqdMI4NDVE6rpGC4UwmKVQXaSXQyRLNYnh9iXq6Lab6jKdA7Pp
BYmOaNQXAFpDkuZFZToUMFVT2CNI4cGHr+O8u4bON4+fDl7GQdbpCKVW8CCPylwl
oRQFbSv8UMWlJ0OBY2YsWM03IYdmnnpkGKH8+JYnhJjAkTTyw4zkIcqDRGg1lIIo
00Q9Bpj07vrJP8b9TGxO/0paOuM2VrWXYXIKrsB+LYkjpUvMF0MgXa/hzBI0X9JX
/yBAAVu96DKd4jLOv3LYLvnR3TIRv/BV3HXClUP8XYeDaDJ4o142E7HUa/DVrg5M
wbi4noavZVv1wo0oQwcBAh6QYz2y6pc1FyFtxjvlCTlPDrP1OKRpPe4Cf81nIsFm
mZZFDEzEANwZPTUHNaGGO0gpjb6fNUVlKffpr7ZTpeuKH6SIq6FVUIX7bWcu63P+
vsVN+xVZLhHQP5kB4LgMK3TFORTP5qMABt9AhoB/7OEsKk4Za+iJc/L54lQQwjDp
JdKzhAOp/K6D0YKFvWLResbtx7hTM9tx7N7yRaH+FLlbV2j/bRp8v/KGCeuGyM4v
tjZHajbFud1W6qmHnEfk9RbT/CfzFqpTwLeEogDl/VhPhhgDzHGWq7Ls1weaRKIN
36gHqkclTTuE6X50Svxi0LDjr/uRYKakSYot4QPwCDHWuSW9ZNQmMhYbz7veB9KI
PndpKAsEgVOMir9UAoD4mIL939hZHVUYoisXTbXikdHJqMvbnZG3L7v2rs9IbvGA
78mzu2jFuSH7ItSF7pRV/ZMH05ehM5cAtVizMmoB3IZsOKht2MHGPpjxfsdkU9Ht
9gJ+IoK6D9fPLhlZItdghafFhReiUKLiFXyD8cpAWvqWeCOhWHuBBk+sCdW5rFpR
vIkALYqR6TfGpiYHZYC7vvFzV3kJBoZu4PJ4YIavOLZouOQv64+VRbrD1BVR7tjB
lV9x1mjuXKyoKSq6D1btQbBTFj+zgLEixnM5qA+hRVXn4kNa3bMthwjg2v9UOBq4
gAsDaX14yqrh977bQ6EyU5iyPYPRyMCxaR2XueWg+tLC7Lb23N0L2X1J8NbeR/qL
HQgxNou0Tb6yGCuk/EG8+WJP8EDbXzKoaP/PR3YcOdvKjzDmryBaXvXj0D+AKepm
vU/luSpjaT3GWMFvvNMYEuc8KT61Ze8HGUZokuqL4FGfQMNyWLp7qX7oAKd7U77c
s1pdN4AKXvsFdcHnLWb4+Rfng3WT6N5cijNanM56pAScYs+nq52LgEhFboVHtHu/
mWQMmOlYZXsV3fMcJ+1Qkb4btRrcQF+eT4ZZ+7BwUybcmeUb5Nqd3m74weOUNjIT
RMnaahBmIt7agXGBQuVgnnB6qGj+QLyxCUZPc+TVGji6R11XVkiu1EM8pjgVxua7
0ZjWRnQKASBPbV5XUQb2jvTZkIEnDbZBWMoJPYCp3OvR748aRWiZ6Kss4MB9rP9z
iUvzP/RWvdYRidII794eW+khnMYY/7DzfDVTE0JXCmwaQBO4ddE3t3rANTz4226b
PBjJULgDIKaUm51NGnnlYC/ssgCmIfSPTyHMkTqEEgOGqRcd8TW5b0LA9z3sr6cf
+Brq79j9dUsow5RUw22x12YhD77ughabdIIy7fNb3r6kyIzwyBJDoyKFaMBepob9
bz7hrwdpXSbIv+RGgvu43nTxIPX9dR6olNsp3vbAfDCVkztQTCZRFbeCwRsQ1Gm2
saT+LPpslTi3QFzHBd8UY8yNuqb+3asMvOdDSSOxboPr2yP8dZBUhqgwi/R5zA3k
/w0yf/bPaHgaKuXgucSbn9l5YLGS1QHYWQ9Nwv9e8k5d3HpUsU+sG1dQaojdhoBj
7zsh22UWO32rRKX299o/c00uOktQWQCSVTC1aqvNoKcek1DPILxYATbNS2XXxEfx
kSSu1TPXzlcWxI3fQ7euiGq7l6HaAmQz7P2232oBFbI0I+m9til2JrJtvg73YpOh
PXzVc509ebnvTKOmQ5stWeLnan5Xmm8mbx7MZQeGrRnrLuSgM1iv4hoYvhw9Am3F
oqThwZ7mGEMklvWVLaJXVdddLK41E+DFNH9d1dH9zXiBOQ0FLOMGKoEFusk53zkh
jDaAE4PUVRYP+nyjiMgEZTUjTf7j4fUIi4Pi3Gau+0J+CKNlyd2e7mY2EgA9aEyx
OnnP1fqjKXXrf7NrG3AzAV2/IRrpDZO4Gj67vDqfLT8Z9w0UiDW5VdUptGNqGbb2
/XK3kQXTa1RYv1IxojQ3sGRn/2D3x5PhTLFeSL7wIizVOhGE+bp4mkjpaRhE3utw
9a0a7zgQP26ykFh7fxTWVRmExNV86ECPpfH/GPghULZ+eQ3RSZzy6H4AUWwQToVz
NDTJmiMOM9u4ZncPVy2MRk+rI2NkYOsb9amtKsRl+kR/nfRg88RPAjA141XM5zko
NTIHSXWAVtmvydjFpO7wpN3yQkpYmRwZh0dtQl204SYBJ4Eh2bxB7SdP8OIyRnHI
zfTT+S8nvOf43s6IYy1qewDk5h9Od8K6ZhkMvTx05La4h/vd9sZ2hwmxhL+KQzHE
EMUU2uDGWyLeQErP0BVkGHAkxLYeXJKHpX5MyrgXG0DCnx7wQMkRFgGE00cVDtVz
gXU6ZwgzQqIGOelLZ3Y5OKMwCbE50Cozr1xJe8fDAFEk1u6wH4k5Xm+foM9RZU0o
BMjx/8rf0089g9CdYIrbcVnmpbhXFVATAicE0WJwqUNrt2WxtUqCVl3rfOslKI5z
TOu9tZE0VGTjboKdWff5+2HB5aDcjDSn55TERUm/Qc7zkFLcndL6bciaBRqd1ZIi
7xf/WXs/yLHBCT6ibsQCpj8Z6H63xOy9Rg8cEISFN8zHFIlmTtGxV/V01oo7j5ph
rMNfeuJEIUk3kST6D7vLPnFY10vMFSNJdSm+7GZaoYo8ipXbwRlmAkDnETnaxxru
oOw7usxzd9rBZiJ/IU4EQWCwxDWnfb7qBZjv+DfCWpLAX/P78oTU/+qNbVSHUKhw
MEMWHBNmV36ToMtYkk5LZ8zJmMKNi3IZZTNOPay1vI/hVdIaqcC0wYM+AbAKDfRH
lKJiRp86CrTOOG+Dy5+cIULvE8VI0fL00Nt0SEh3mc/MT8uHV7pkxVgl59viR0gJ
KA/pUnJCfnPJstZLDz5nXTgcPuZkX9VhZF3fY71Q8EBHnNqe50m/kw9FaNjfTJIa
d3bjl+O4jMldis9OlZWcJiKRlG8kcktOFCgdxO9V0D/MMBXwOh/X+HlvtFpP1mXv
uua5ipzmHyFT7v9unZqcbSq63Isw/km2baC7WoctoV8MvIhei0u3/w9dNq8prXrh
KfTpFFqybjW4Ga94P6fBvc4D8gQQr+q8kV16ClYT5HzF/g4oKIT/u38EkhkeSPvr
0e3ArmE1TvMy2nKwKgx6g+17iZmvw6ijNKg/lfKEQEb9PLCTZ/+nUkAPvKbfx+MM
eTzNWSt+ghbb9OR4ndGp59/7oZaOAPBGjkpOZM1MEcSsq+SphLzbiYLNCdXLjWsn
ISdGCsSs8SPBVNlm6oVlN4jbOO6D2cWzzZMl872UBuQXVmuXGtp+RJHUe3tmmQnX
dONEkeNygWn+gV0DVXqnojEjF2K47KbdxkwB/NQOfPNrns4MCH0d77CtneMruVXS
1U8+KdNyKZrtXRVL4YnpEKHHPAl9B9WpKHxYi3VUe3OXG5lVRmfwdjztXqHOJM8f
abrIvxXDoFmssMU/yYthWjnqSujhx266irjI8c7cdWtmQkpIdYXGJ7/IPUjDbjBm
5X0JiNajn/ovhu2aFkLaOPzP7fdXskp1mDhEGP/B0FVPqu7k5q2ZUXYc8hIbdQ6g
c2PvN0nvKA1hznzEF/ntx9yAGGaXurtwn7lvzty547nr2ve8lHdCyA0680Pfyfvl
3vkxfXN1ncl7fICr9c4Lo4YB8rDv62Wrc2kjlY3E1BI1a3BpcdY+NPWFaktYCAV8
nHmprfnTRzAKKXH+FEUBQQIzKWrAcTZ8cMj4AvwyxIqK2A41yH+w8pDrLCnahSMs
vaaECJqKEhxQNqQnKgoPrhOUaBDE+myGxnPDDFkthSBO8vv3L5ZdNt6ai5IWBD1N
IOosyro1YbYHENPDBJqfocbiQ/CvraNXpQS5jR9QGwLB9uOZ4Tl56HX4PkmWXT53
P7vSpAK0Qt1jjyjLH9jlI+boxz7Mps+ieQWS+MscmdbPoKovO1wzAakJiXe4WKtA
ExJm4ym33uH9gOMyh9GGxPdUzraJf3DaFniZLM9I3c3Ztv3ar9e3D+oPLcuo4qxG
kVsfYId6hiK5z92T+M5/EjTuixXeyhqmhIU1Bv2SLriFo9Ohs4+wiJBXQSC+2Yyk
jsmGNOgJ8R5fuYDS4JCDaJrRKOBcCi4FivQXa4gnYZEsE8jjqeLiMxC6Xg9lC/Jz
bgZ051F8orbfY2bgeNCKh18Jp3kRDMTKtyq1P5EQAjL4CdVuMwrhUCqXryNhzmp8
cDkHJ4+OoGKAlMEAOA69avFM095p9u1fQMsvbnvFnpyam1dUN/XWtfuVG6GslEpu
sQ6RyzKGPn9oPSSev8TcDvsRAi3RH87LuROUN5/x0wC4eJmxgGiHd6tsMFKPH9YB
Ir5lAQ9AMdmegbWW8OVmfEQg8T/qWzpi/EtQrAvibzZozm2i0msdnG9gjAIBrCqV
PowYp6F6TP/iwJUm8hmKpqjEZltfHFxZjSrsrLgeXL0Z5lzndXcuaf2+IaIS4T/T
H2oLVYmtLmaSx0QazLXDID7tfX0imk9DI3fsq3wvzH957dcibZUd+dFQruEwy4/n
W1AS+/UK847OWnHc7yehPJ6d0bdJtXpd1+riwwcstM8lCkP6+Ge86G5t4NUIK1og
B1OhFigbWXFfJQspXDebQ2Y6nPxRZ3nPZgDfuZ/V4v6n8FuUcp8VMYAbLIFEXqsB
XwJ9wZXQ9hivBQmyfI0ma2THF8fKmA32vlusd4bxNqCdWObq80CyFJqfmh7jeqqS
vcdO8UDQrzpTnsXh7Z0Wh7VcIQ5+3VJ59WQNfCYmhlnIrSoPOzFhUTo0x+ZPBPXe
V6eYibk1BGzb2V98I/wNgfBkpjyjblMoNHlUlKkcf29IujP2HavwJNRgUx9cEWB6
0pZmcWHGpIEds9RgKI3YE9+dLzj3WChyvU4W/4ezqtMu/abjq4NmIAtNeQ6q6zMb
xmVBz6xKHjBbZ57gYs+ytj/S6X9hD8NMSbapJFQ7CYf54xx4oKvfqDK4B5bL6/qr
Xw+YGyV3ryLHJZOmjLXATQavcm+WIK5L9v649PusnSLXpuD65siwi3VntD9CVpDN
tVpFvH1+cAsapz+9NwEphUxpgvOVX8HPNr/IKxq7eB8v850w75uBPQMeO455lsEn
s0izyaQ+PiepiI44qOQRjr8QoHjyPmCP+8Z35uEfPe125Vo6amZChG6Hz/0PKLQX
Xn1VeehDchQkBxwGTpelAXVev0sm8oD+xs2ohpRAM5oxwPmjEDSBWrXuC2M3LtVf
7ALRO/CpXtCNaw9h+UoD0rLYSYo1q/qQsYhFxW13aek2Ki0b7WEnCL2773/+yvzh
/s/W98N7yZXM42gOIcsdNNvRAk7BUZjNka9UEXAMrjoUoQxauC+yO9AepAvJQPbP
TT00WGh17HhxGyu4Ja8RhwOEUG4IiGA72ESD5dEk6oAbp3LGmqmjcKNPSAJZnu40
FZm8NzgrZAyC9Xaqvt8mf/4CbtXdlfV5aEdRayFDW8iQS/ttOALL+O22TeFCRtmz
EkQgbRSEEVpVKk08zBq3eOYe+Nt/MpuXkMVPeGe2NzhuD7PhzVHWf2KA4//Nw+O3
TLly58eU7O4DnJo4EbTN0pCsuWc0+HrUxB9SUZu42t+x55hSKF7Bc+rS+4Xzmkkh
IA8+lkK+gsbdup+Ts3LhOSdqZiol1/m7Y/XM+CMrPRaWueFPLeONX7FY9smOwD6+
5wSK25IYQODehVZ8KHU4oQymxKxBxjvfffrq3GtB7MK+jq7EzGs87s3++z0W/jqs
jS29Hljk63l/GEhv1/dx//hMantsBP2j6KAS9SGaiexhLKXgkaeCYL1Av2RYLIEn
86JYN1z7CLzTpVcYUP9jf71aJwGYB+LmHyveUvWUtrgBHDLVi4k+3jFEosJcYoIP
7gxVA1HxJYzRWZd54jPg+SnBy4dVmlKOHIkfSSmTkoXRDjbdzX8lWsqIOMWxH2L5
0IjGzc5U0+1S5Rrek2VJu90/56sOcQo12zsJFC0PCFE7h2UrrLuqcIcdCnM2QP9k
NGVUogkpjdhfgWhk+i/u5NoYhKMzHXYyY9GfSPFH+QaqxJOuP5hq7hM52fMXbceK
5qHfi08ZhSRlnQhwPIBGmfR/QwQkxFZAkY5RXq0dONbHGo92YBgmvB0+Kojh93f5
O07pXK9EShjek6Iw/saYTWxujU5iSydiGpYoMkJuG8G4UI0dFpkJFST7cbiZOIs1
LSSAgxBV9m2a9eFliKST2cVY31ij6Upy05c2HqLUQKar0zdH8MWQlwaAJqPAaRQT
Fdon/3GyMZHEtlOWzpPhpgO1NvHgk74phnZsGQA5fWbzYi1tzRg1OqOt+xwrX5rk
fRC04McNBG2tIpFpdIWxzmaw3lRmoubQ80bTN2vpVk+MSL7Aco9ITfp+Hmc08lwa
JSKl01r2wQWv109/RrUoxb8zVwI9qXL1zdKWvL7xWxIwuHsgwYotH4TNJwkh8NXw
kWdam6yYk58CiD8BpLFjiMV0fVdwbVuHGWkMS56KSPjO5AoDSaUX3oQfd3ruO563
4C6XldAMQIiZDS+PfpkPFMnJyv8URVdeoPBFTK3H4khQuzjbRQwyZ+MqKvrwZOpw
Apdig+vBEnnJcLsMUUwpillTET3Fn7G/3dISJTFwMyE7XswCATkSoyzJheghEgeK
lYYgS2+9ZnjGOyCd/Wgwt2vA8KcmZOKUQFvjjLNuc40gKA5nk159PhvHyhoSocfi
l1aQqsNW2Hv8T1TyjzosU4TUkUi7e3S5ELnJaMHaF/MYDp0MuevMy7uk5w9WUuC8
C2uATL6GZ2OFlkGuE5+MaaFZwNccH1/HQxHAt+VCYhy4Nu7MIVHPFCKSao05HUE4
FcfUT1aXmh/c5Ic1wJd9Eib4fLy8Baz+96wayWuYuzmrCDbLFos3HQ3dN0g+ToCk
aIvvPnWhHT+1sAS/M5HgOBVTZNzpgrIbAF8lO2j5mviMb0ny0QcUA1ylFL1GPoA8
6HiWZ41npj41rCMkP8u2fqXulC50GC+TdgnjOx7WvE4LiDWuwHDsdhPcOTWnaAJZ
TVVipgZ0cFZxO7pwg8rPdimM7UFPstx+7w6UFoMIFYJW7u+7oJfHxKrLZLOThFEh
eVeErpdxyKgvaNgI5owCNXJFWuIFTCPRSY4dSb+44BqMmBbqJfPZYjTcGkUME6aK
uNmULjIGJPjHTfko9uWDvNRbcpmzQP09Mwqy7RpJPzfpmrxyr+6Pqp3uhp8xkUaX
alM4o148uA/7FrQgVPA/PJF8SEXPwny8eVJD3niVZujLOx5kdxoCAAA5TyePlVSx
XSjF9uZsdtkXN/O55CuVnIzbvniFhm9FOeuVpBoz+Os17umcEgZb12c3hu+uK+OU
JBzsvN2em1mLis2qvx3xwLPkSluWN+Fzhcao5PLIbub7vD5bIRQFMjvHfV+JOmgT
VjBlfFLPUMtGzjzZUdLaF0gYtKrO5xEvtMw+cUdvK6bvi3xLNge8565mrtfwc054
NCAEQ8fdQAitP+xrloUGZX+5q6DSWa9nYldQWeLV398yvMYdwSjV8Vr5aGfcNMte
KC9q5u/9IreDwAfTfkJZEX7qo3TXN28iOVCW2Vrywt/TclX4BpOpE9xLT27jYGsS
omQlJ7a3O3GCM0K/RjOtBIfRSoNsWKqW3SzJKvZKyXxVIQ1JA5zl1F/tJAUkClCw
dzkdykKDpaD/SVqTq47r0HarhLZCb+U9t1Tdj8dTwMMp/Yq35bsdTdBJDJjfNtRc
0C3Szqx7Oat4JBeSURi/xt/3uQfQgJ4Q8BIVYDMBdL1R5lBs8PYFHMvDAGROcybX
momA892NFwk7UxayHhcsE+hY9HkgEj20UZGzq8QnR31sc3AOG3FgJWf8nxCWPFrD
PbHKr24NZ+kkY0fFQ+943Tfdg1VS7FK85Gb/gYN6UReMbDxBPI4RVW3RSmoYhFWg
7CpjXE2HxIu3ubtR4vPYo8bQJ31P9EsDY/z63XY3bvIsskU68xOv2fbmlwJlKUmM
wBcGAg2eYFNwOykhjkEtg1cuxbmsBQ98zutKI5aGCPSq1gW0ZkiodKJf2MRdYS5z
HWlfH9XpMxxOQ9ZCU5fwJYXup1OctROGxnl6kmOx/QmmCGfrh6ZfNrcmxmHmWYpF
Jg6s8zvjMdLMGhhcFNMyor1sh+IG9MPz5dW/WBy+APOo4G5ujBckuGyRPD8VONai
3qke1KMSZMxWoJIfRXJMysvvt66e8xx2Z67//pXdCsdp7qf/Ke25kjsHfTsKIHm1
YM+MU3X3u0PX0wVYi7ag/NNCMEbIExdNZhUtCM+QMiFKmKzbr5e76065AGuAS8mS
TnZrBMiRPAo0E6vrDBLWHLghSOPDsN+nJFlbKluSRqHArE/UwDN4xgSHguoRo2J0
2rBT19nx7rbLGST/lPSCgB2wh8jrakfy6+glWnYWUQdIe3Zpbx40diBUWzlN9/q3
tbv2dnlefT9/X8JAS3gyr/psfTpkCi4cxJzmijFwBkbUn9Q3Hp4Ki42EceJ6sqlM
25L0rKS2rputpEn0l0lTNmbPePDK+D743PuXTAuaQPaGuDPg8SC/xT3UzNWQk9xm
1xzs7LbxtPu/C5e4+1PCTru9RauF0yjicRR6VPl1q4UdWnCKMPRmvosYCFyKBmf/
h3K8xL/jOI92f0OWW5X9ZQ7elQz9YkkQDic3iKXWihTvOla0biF/L6m8b688y+L2
hH/di2/TZUniI/PbXRGVVpbHPxQDNCnzA7l3AQrVUNUM2ozOe3Sjn+GUA6hNNGI2
IwODBkUbViBR5GJ2h1mEu9FEvTh+rp9qmvcp3pRC77Op5p7Kgwx/HifDhZ1vPaCe
/2dcyJ7hveXjXgSYUYOGO0oTHzy8AB1acm2FUxH7jTr/UUg7Vag81VxtxQYfUCgK
WqHMGaoqivsZjmCf0izJ78AzQ011/EVXD4J3ZxINJPDJg+f/3x4YYdiLW3I/NvuC
Phatt4SpQbffM8/GHhb114MXpGSzw/3b6eMtkGibo+pRX+JxcIOpR0pc0Ntlc32f
HQvLbBODqsly307sReOLMqCb0XHxIzZ0CbWt9WYkUMVH0LgpyzwJxUdJZjqBEWZM
Lo07CfkHoieBb7pXiw8OYs4QRvsZ530bi481XwPOdL5BTd5vG6Gdo5dARDuI/93J
3mU9XnZ7wtwW9UjYMZjwpHl7RRMJs5GcXxNvRbN0aiL1FiWPEPD0+qzDAszG21UH
iKaeR8ygJmSqHrD2X34O7tV12llzZGdjhTgPgQCmv0t+SruE1YhlHg2/+LSik7Vs
T+BMRK63maq2Q+W4nqB0ci/ULBKKRiicWEp3wNexm0eUhqrb6647/tKmBeydkvqZ
w+CgBgVEspKBrjQT3uuUkW8YRxs8gDGbBOexLBFlN+uK4B05y6kfkAp0GawnErLF
5Q7KJ8j475fa1KWyNVQxrw+Jn2Co397n8B4Gdb99HZadW+nXYJ5V9KJgD3kjsmv0
hw+EK261T8bQK6TFQfSat5SNXLv0Jkm4vvn6thJzNIPrK8rgZsvPohj4qfIStWW3
KU3+vtCQQ5VDPoGFpUOx8epbXrgHkpQ6EhICeKuAsejTRgYDhIM2cMTbczYVeAAs
P7NJV1xCbuookQoG+6iCjx5ZmpRagsso1lqV3YO/cN8WuibQ3OZaGDtbZt3Oe0dk
5gOhT18hO9385LwbeINuAFxgEUKqAaM+my8mtng8A0Jb3NZ/C/hIT7+HKvIKOcL9
hSyegX+AKe1xT3SrQ9ApFR8Z44LLT6SdXUdwPcxeLjaObBaSvVLdydIwS8dGFw7q
oUJe2yZW1wGBR20Jw22KGkl0W1+1OCDmhYn8DGchkaEiF92khIqTw78pYLzOK4IB
2zAmmiZ4DcyInk+TIYn2De0J5d4boAIOz84sYxUmRRwpgacV7t5vUf2tXRTEeT8X
DjZWJi3nNYQKhy6/w9N93WiNfxiNQX+DfgwMzG4WexFlBSkJNU0KVttzPlbSKROw
6mfl/bQO9WzNmRv/9L7aLfNiH0PE0W59H1wroVFMX7hv/Ed6EEGSpwmXkHAscEgc
7zRrA0AyZa+s48owFZ1AVmlqcvCiHyVLjaNP3222hQk4eZRQ3A/gt+qDNCaJIy8l
gdzYRF33q+r3H8gx8H7rWPxg6MldHiLHwseaF5F1htbCnMl1ry/SkPKMwkg9mNPF
1XwRkqqYfrCyY8dleiEGamtwl4wZGZ6kFAT6PL2ymmG/zrLdRFjzv1hyIPHHKv80
yXBwjxOmUXi6pPE3FxSRdJcHC5UQh65+LhPJZCVB/w84ZTDtjhTDQ75GCqIlD54/
jYE3M40ypztmdsthg5l4e0bbo9KZiM6nxKndjHo/l/s5SvOj8T/SoWKAPNOqviaw
By7u7/Ed4uZzz3RXEiBqd+RAj7rOYfPf+0wVObPGDEgx2L64hOiRJucLZeUVFNtn
Ib3Bg8GFglUbSsefntLxn+4zXLmq0BRANgoT0lgUzkR2SAE+iw+5cvxU5xaZvIGY
d6Fyxlwj1cT9ZVDNnvAnYqbsRZTreDvtu0J10AsDHA6BJguWmVbWj+qsNSDzMAeV
ZOWOsimSUQX9gexrs5lew3HbirBHQXVzWnw0tqt91Vrh3mQir0CdAcL1TpgdlJjo
l2DB16Clm7FbDtz+QXJN9WbgT4EzzJuz0fQthaq1pV9kNsbR6Hh1HHWawDYnsion
t030pw4E5pSNSjZhAYXGHC11nud2rjQ8CYcyl+83uv0dYsEsWGT8ofWlUKUCWgsS
NFOI9b2L/DMVf+9PNgJdPsfnDCJG4py5WJTErj38PV5frO7tUjrAW6Vkntu2qyuO
25bSVA4vnOB92i7SmjSQUSqZ6x+F9O3PgkxF0E6Mtq/G5bDxW5Nm8SGX/4rvnLlO
aFkvLVNymJzhN+PifgZExzlmj/lXbfpRx+oTU3LwfVvPliCakoHamZJkWkCn1TtX
mJd5WN3j5tks+TOlOhsdzf2QtcBCHmAoNL0Lzc/eWp+zJfEjKYMjOfRG7ANdn2wk
LOAe2+/Nb36e7HtXaILZwXAFSHeL9/aQsmaCIGvqm5ies2HGjzbSq00Q48FO3qLj
XkWRihaad5sS4Iw1h5MBDImv/p0Z4Enwvk79pWo+URjybsJEyJItoalrlvxQ0cjp
OkA/6XW3FcZUv4XaRHkYhfaAThkEY723srDRI7UKrxpYGMPn3UNsZ/cOLfoMpwQR
SPgyY64bEdZ91zJQU3kRF6xE0JcAiOuiy3U+7Q0/yEkWm461aKCAsw7FULhOmgta
Yy7BQfju+GlYzxAbeoDyf1p+FD2b53j0nwNXyjO8B2/XZdVBQQlbbgrSs1ikcDoS
oFu2rvLogX5KX890hWOIbBIcCbaOab84peCoHOGn5ZL9/IkOiKk5tl9vimcUKs3W
jZTakhxL5iuvkFFG42kwVX38eIO68xQBKGQqLziptcy73Nt7N2NyAzMdhTfwxeih
eqb/HzEVxWWMqaWiCENK/8jqjyk7kc0o/hGADw+VJD7AE2rAIDodzpo2In1X3im7
6o3okM+1zVBnW+8UjyYrLM6CTsnEYrk71qkqU3dMwhIujpsspMrrBBN+Z8Ww88ND
h0xJONNEGN5ZO3kwq+6lr9DAntGtn9ZTUCv9bhMU83TS0R+GNZkbh8+16d9IkHc8
0hl14HFBS0DOeMjCTZZLsqXYNFeuxZWDJu8XJmLj8SpItN4Tj4obPKmgvW28sCjv
CTBnEQfIY25nyFKlJ2+vwuw/2ztHcoiR9QuR7gKG3M2ksA/1xOgd+4u0qgitgHnw
P9/HOctvQoagiPQH1RXzI5gFaqP8Nlz0KovjYycx7t80TAT9/iHcH3VKwt1inFMr
dFL+DWFEJndafR35Z1egRWdYkoHxzpq77Vf8YDcQFL+4Pn+r5eDSnYtDEmY9L1dJ
Uv7f2yioAp82KRbehuP56uAq2KRCPYqEF+tkXUadGjSDoySdWRz5zKYnB2jD4B2r
KQwq/7ggrrMlhPmdKmXwzrnTjBNIkhWwltl2oQ9/+MnLAX9+ZgMj+o9PTf1ZP7nr
wx7i1LwqaYinUwT25vkEBxLQVSgLraBMlw83EXZr0SOf8h0cEuQAKJOFP3yc/vlC
Gv/nHAPQOYc0z9RnYYzdCGyqOZe1EToiFEmj/a3Q5Pkl5cEEymGBeRQTxK7wk01Y
YgpfTWckhQxuJgtHhqafNHzL1XOnSOZfbzsOKMow2iChh38ZtSeWhtkXjuauYsAo
RsWI4Y6psufpqMb7ChgXcU0cbghH8nK5AoIi7ecetWV7ZoOqXkJWd4HqugmL4Mif
RIlP/voX9JZdihGhSnpx+e5wt/zZlCYdmjKzAHgZNRj+fXr+bM1wloPxewQQgSaM
CTgzmXcG0DXMKACcJSXN02Luc5uEHZ2diopa1qXjfaIUFacx3zRKdrhDzFOyMbEl
R2hde7wGBwGAXB0/lnKZNa/BeGRxDcPBnP3SYM4HvqHklHLAL8ww+D2FIdRQL7xk
z5NHN8MeN+ztzF0amVKZYPUJcnaGR7PKozBgHjybmCSzOEun3UzgS3vGd9+Z7f7H
lhnEQ5eDch+0EmyAD6NW6rCp1j7uplOdazOT1hScyYUqimszpnsF/44F95En7y3i
TePqXcdyWKcBCORDIl+LqYPFZ6a7jLrDWehPZB8cqzroE7qt9vSBb191u/xi0o31
j8QVqT7HbERJIWsoe9B6ubQWL8oka9fDjGJoV4H4R50noq0cQbF0S89U5I5YHnHO
HlMJjizU70gVbBlU2vAfu6AanKaiGhnlutMlL1CTzd3JAYOx2+ENqVR/ch6sQC1d
WdeQ/cwyuBlwQI1oorxdwTe4Gb6DZgEoGCc54d0fdMY8+RNcIpKd1f4dkIIwlD92
Dq7NRh8dpweytvGaF2PuNezX8R9D4ZQIe2GsbQ2CiQGPCXEe008divXGUvhBQoy3
IFYCJIavdi//3JoTlkQ1FKtvdAQcNqMlxS6/e23D3DE9nJTbsoIkaF/MfjxWeK3L
ZNqW/4KSXiDfMBtOYzVo0roe5+B6Z+FuZUq0d/d1dKZxDfnVrR0+uHQbuIBnxTeP
qq0HsJwgspBYImPw4HyUryfsGw3rXq5b2M8sherwB82cDJa+Vg02gXh3MQpnMJkU
QUy6z08xJuRzrPCXvVzny7PLKIsSYf3J4X7YHrPTJZlxHW69UmYLoimzVlfZE+ud
o2ytxeV0QVIwUidOW+FJ6r8N5vXD8LeU70l20OpbTRZDLKHYWWfaY8jBi+z2yCLi
zl9gIrhbfZ8Mxa9r7cAhTr+ID8Gh/QMolvT6VoRp2T44hSoiPWzdCM5qXN3KRm5J
2MJ6OfpVLA8fSRxXVQWD99tZRB83usF+LMapUDe8O9ZqduHaNwqv1cryIpIxNb5z
CQoOxpb4h3gxqpfNzdb9cTK4pWlpGI/l1dCkUSNvgudYbV9PrzdcFxaE6LHf+8y/
GqBhHb52+wJPeIzCITPsESqpzvsTEz4/nseXMU593V9qExHcNHO8CNIiXu/MLj/3
+0KFGcJOzxP+QVLOcfAz+Iahl/+1yjYNtkroR7Tm1+DmG+xSa3ubFq6+s4mMFitP
qMu6rBybz3Uv/t6hhpPytfOal+0JmEK5MXMkvR01zs49UIiXxgZmTneUSK0uph4h
zkrj/RMsIEVXP/4doudJKjjhb/EbZRbKFAqTqejKJRi/kse0cfGAB+1JzcTlOKTv
TFSRezDXgiVw6V2ct8+XwKN++tQj/ABqAICp+fqbyE4il1reufsTuPPB3xuufakC
OpsvBDQ1FXesn8MjDcY7VPBDsXb726OaDoOp4lNBAeh6fGNfE7BrYvaz5aCFbvGb
ySAGdvYheuFIN30L73fVbEMiKnHuXwZCLshKfTC60odux5EDpx2BUmTnRhi0osCH
6kiPlSPQcYc6Djf6GYWyrtuCDA3WDoXikh6qhLBjoscofoXXEQcMPMuWUi2Hgb/t
h6woIRhjJYX1KohS4tLLtJ7oOKhvT7/50iNPjgXhg4ZG2CCSuXuXeybXHgnGypzP
361zADw3tIRSngewyp/WCAtplxV4OakcW1RlVVCGWqaYCFSVpF35OhGT2ArDiJd4
yZmgFIR5zD0DExJoeQHZRHqT0dEKsAOTBD2sZwPDXu57w/zCUaTNHqc4a5lwlURD
o8yj9ENkw8AWCp6XZjmlcDj5l9N+iLCylbCwEC7PCufT4VVLsb8BKf93xBE38Tl9
/EXrA6YLwcgUvp//KNfhqX/qJuAQzXnwVfIZP6H4LV2+Xjsqc80DZsMaCKAtkkAv
vV9qX3hXFmulc9rE6gu8qwaibpSHxYl4TPliMvrjRecGCQ6zExEU+Q8WzaPIxCWb
krpXu2YkANRoaBf05GaLItgM2eCipUQ5ykLrHU5ODitoORTyzSQoPHkjNpLI8jCR
d05N2A071qC6fhZHXNkspfsK/RRz1WECw/gvo7mfhBzDYar8dBd6IBUBZ1XIA4j8
9/tUGM/+68OQojdj60eEXcDOKyhekedw2lZ8azaj1j4CTdUm8O6F/ITqhY3gUqcF
5qFdF1dQOI9bC0mR+5OkOBXHJMgi8ynluTQmBG+A0Jof3l7taROZ3OoZdnNRXBRG
XtQOgUQgI9YYQNyMLlL0FrXsfFchfQ93Uk+nbEErbRGuVBwvTYKD15SJWMKLB4Ju
tklICvIBjh8D8mntzoMuEhGSgW0+K/a9hpTSWopcPGtQo+Hcg7BbPg2CX/rC67k1
CTr+3lBMQ2IFD1CfhyUBnCu9mWa81eYOfedvKQQN29Hxf94zRTZUwKo+wG3+1yLJ
n0eWEI6bitMGlYs1OkV/QDb3Odebd4m6/XVEuIRPUEDtpVdc3Df1KhNuuMf6tNaM
E1gU9Zi9fSGEowKGAa8znDnbmwvocjy9auXxvhemncRKqGe/H792gTWLLckSzDoX
vHfbedAg2KZANUyaNo5PGigjDXKKd9k/fuEh9Fpw2ZqS+0OuTmgcpbcf6zv/R276
yToxXENwZAD9A5OtwC5tDK1wnTvaFXqNay38ptnTNWOoSQEF+VJySeGaiZ3uLWwn
dylsbKKQ7OmTgvgQGlPKyFpeyC6MXq/0uJpDTlFwDueVZnqvYWUFVJ7rAg1ZgoiN
h7JctZGafBqsWWsWOQE72uRF+wrPkpZ0hXpg//k3cQwsTuAJ7X/HUuQS1KuR2ju5
j55sGEuINc2vTL79fMKKVH4yz9Psytbtz7UcmQtqqWUccgIc3y5IOAz8343f8Qbx
LtiiHfSmUnkQYeI5uPZqufUCtD3wsNrvTtoYN5SchiafWUzKBoR8azQe4Rm37YbP
aKFkyaCpYIoNPfdPeg+vCV+EgArH8pED/mXoyVFNOqBev6gVQvPhK3gmmnMHbYYW
VDz86PRsJmMsR8LvSZuRpXci8hY05v5um2ebuNLm8ienxwZhnolvfGiOs6vA4XkQ
9sDNzlt4pBHWXq7Bvtp67SEfN6bOvG6bsNwXQ20IvwuT6OAwjWT2JzWr1llApI4k
A0REO9HTs1HAXi+WLw0/JXP9nxTWX0Pz/j4hhoUNbdGRm63gkV3JBsx0WoyDMS6t
snKoGl9mncqCzoGXvxyVWbpIhqBTsV4SA+SM4ZAPTP48MSEtc8yZsu8qKqlLHE91
hM18NhinSKhEV9K6PWOQ/DoeEOdTj+QBP+ZGuOROT11xjwJHdrotVLaxB4NCuRHq
4YY3KEh1vuq9PRrDptorUB4wu4et0852rGuuHOw1kpp/A3i/+OGPs0tZv2AwRvmk
gjRrssmzCQY8jWBB1RiaCobWh3uluxCcFrRyCZIfeqD74q/1iP7yQxq8G7/M1Igb
BSVtwZNqsL08xE1OPO4WsIgadkclPCGOEs6uxad+uqpKm9TugNXMNrMcrl3BkxLm
2Mqqc324E/IxASq6ECNg3YYA3P9m3Hfh0gh6FjF21rxN8yDBsTWRCalXpE0AWXq4
DF0afx9dEPlB+FATGuR658pz+sTZRKbmAXC/2Kxj0eytATJGCZobN7wyIOeViW+u
WCxrtFc83hazG6I66zJfK4arTHk8gdQsoiA+2KmLyu2um+AetgJ8GWY3e2rom1e3
WYsTCfrZ0c+0EylMxZiJDA06LdCbhuuVJw4x85Vjh6xcdLlm+Sr1hPaKH6S/fiMo
91aCQFesyWNJpP43x2LZglKA9SYxHaEtEXQzG+BVG/mOw7QdCCd71kdYF3sswG2q
thZwzNmBWpn2A1OxP16lbw7q17MfaPzTi99TnYtcFR91yeeTs+QHflSZKnyfbYs0
u2dZrisMPYentRlfppndskoktV2nANmd6hIi72qE6bZ+lTLPedYSfgSeNO1GSDAc
QKtzU9DvDZXXWt9RfNqLoamb2wEXvgw+ASAKvyQjEytBXT4aVaZ36Z/hjn71RqyU
k3Hq3KQt+Syr2Im6oI/gSHHzutPxpHg+ssNKCdetuRHdfgjWNvbUEcm0X9oMHLS/
Bkw2rrL81whuXmx6swg8tpMwklvB/At0o4PR2GkLwJM/iEQQkeCov3lCUbqZRpoO
OjGqnOCLsnZe68hV7yRKLPeLfOVqyJJlgpfg59eaSSAhHjGEd0portZ8JFAKLo9Y
H8V/WmTKvbFMpTc7hzWQy8lVuPTzTE5lMxIbC4TENVji/O6MXPpnV6Ch+t+NnXsk
PA9ddrBu/YS2I8EcfsC36jAx07UsfR47emjIefVJRR2L36mwpXSIWDGzw/EFz91P
F1BcSfrtky2sPpCnIuOEiyHFM8Cc0lPqBq5vMV/noKwCz1hYGu3f1Kjz84Hdjgh6
wR3p9JLZ/l8A2EQJJW0dDmgziP9ywNs1gRTR/XHjCI3IHSTn5K24x8iRnFuGOUS3
2SMFhoibKr2GMqYJRU4zp8dq6yBiOtGLT9Btd9o/wnUt94u3ekoHs3T+XYcn7acZ
pY6lyTSwimch477TRdjxum7hwYBPL1q9b1GfT1OQAla+WBn5Aa0HbUv+KnoaXnP+
LShpOO/wfY8E49ShxHkT5pf/FcJmP3eMD4TBkEN1xCf5EPWk8QfUe9Q86SVRErKB
ftTrAXMHuJ3pzDwbGOv6ddDiRB5+wFbfH3NxXSh6bXmGxP4iYPB3QiP+8cdJRI3J
9fSlcfk8OHSzHaCS5igt9esh8bJd1bOgqV8JoSUBa/yA0zrQ/BQbg7qE1aQSbB0n
7BEYaKg/QcefywWDWwfZtDzdA8ibK6I4rTqdeYRlSSqRlO795xaohtkpmfdhQmjZ
50iGzQLuh7oPIynnUr32gsEJ+OexUTDcYZKvaORixiHfuChxzkklg1K0QeN79Wm9
YYZtssprruzY1yEaOzXh6J6Cyno5ZiCXjyc5ZuuHC5yZajl1tZhtA/VqBuhvuElb
I9MveZbqAixsyOeLlcjpH+7BvkPpy6y+zU3rbk9LhajjovysHnAmOfKZ/vwbEbEr
tQ9Zsxw1V9emi9uJhib3IEEqaJj2MwuLBgwFFHpvj+ShKm84L6K7zbrAZzs3KDTc
us1/X4PzuhBp02TJ4cSxykRcjsOj+0O1FI50obZqJ8LRFbxEsxSW3ebLF2ijhsK/
hQtD+bcT2WyVhj16nTAggNQ2BYhKB6bPiUGYFOOkRVrjTEJKvdvLb7qFhaJX3FXI
T2p6rtPsefDdIUjxz4hx3/MfFRHmL9H2806l2E6U+iIL/NSmq3LJ2wKzDqn/dwWV
i1gM+9675lrfrePq0ItXdjvxVUqhFkibh2WWGGOt1+0AkwX005YjR0d9qIt1Rmb0
+OgqghM2N8KydaEHfm88jQ8+5h07T2yOkI6D1p/vNhiSTPy0zY2hBrwwvxEI7ZZA
YycWyj0caSLEelBnPa+2+hna1CYPpSP6r51cluyf0B1bQbTjggjumgSm33RoSk+6
SZLEN70PgLmO20sg+egZ00pJEPB/vgudbi8vh11/FEKd2R0b5prBndKzEAKoaP1P
b71KOtYaQD0Z9fsHH7PlgoPrphMro3/z86j4wYrWU/E8Q2DQatGdsjnKjfpSuaLR
mzRNL4WuRYk8ehdYFzm1CarFNXmOlyrDvsi41eJa5a9XHsXIi4RMqqjgFiJigkxN
85fr2nBl1KzhPPURALhXkI8uwLXePeUHA2UevXfin80fgevx3Ixoa4uTF+MWQoT+
mSWTj5RLGb08VzYxlXX9VetwPKjv9FBTxAYuWBJaO7jugmyXpP/X/RwmNScZ3PW4
Ai8ox/u98MQdlB71mLzLctxPgPW92ZS9fKLjqen/qvk6b51B6lXtqO29hJmTHyb7
zGQgQk9y/8PtlVFC2vkE2flnDF1ru5jSHZZzn/ZXolplmzZEbmX06mLmNLsJWycu
D7PEeHORvv+RuBb65ZtH85jx806JWFNic50HVrquWOCK+/eheSoEImQMBsSOI+s1
aWrSohulsaMiU5YNx0jZlH8MJQdZbi93t7vNEr6R2khhzma9VuTu/y0mDs3Hv5ID
HR2RlFPxt6uDlpdCpsM1uY61L4Lj3Jhwgc5NIcHAJm9shaWydMRFObS+dOQ3zSFU
xNL+5iloVofjZJWIOcGXxRz7xWWEKGTOZh6o/LuIX6l5F7POKmDZ2OVu1Icl32JC
Z7GLUDjXY1BtV7j5iBz0pp3pM7YUwTWXhs/0BU8XarD9yxxQrbEEH9csNnLWGgYL
kcInqYaxL0/miqSEccnfoR2C2lmT4rCmVo7rsyare0MVb09t1QPm9QoZ/vaER2Vx
Gl+HNG1oL1TWflPlpf0oLLaZyV0XPW9W/xrKuT1K1T7FSyShF5KzZqgFjMBxj1HZ
6QNbWyjiUzpwnakWUFTeazei2Jcf5gk9d0T6rlBRBNMKHDURq61TXLwNrw+9HfKZ
PppuQD+mAdQU0HgdLHYV5JQIJfIymT4yDJjEDyz+FHEru83LiLSiI3Kmu3887bey
ufr6R5uapI5Uoun2QxHCwF1rld5wf4WmUmbUaB6R6MSo7M05qxY6a9nOrnVpixoi
soExuVvgbM9q/YnLpzhsyD5J4JZ5xjv6GOGXBZ24eo768Ddxhm0T3wrPqq3jDklB
HxzaaTTHq090B/WYQsEAtw8H7ciV/hD7ypECHI4lslVImDsVWh/xdTaLvdnQAEjy
+sr8OrWnY8BvHo4RDniWAk4Hm8UPbqAwHxLZu2jmBGzlhHp4VUxbA/HFrfG15cj0
RhROlLRwT6Z5+57qcIjA78BdTL7kTT9keuUA/RCQeq8H8YTrMWlwzveI4VUvaLwz
WsDgMfRm+uIWA8kvBB/c3dI+vN+GMg8Cqoc6GmA0FsZmi4YjD3pwrauImeyyrbud
WLAeGqZdg3zwngPGShUqyFuRnWKd4u4U9V3qJONZvhO6xflKzDWIBbUCcii/npHX
tvY9tGGsYYYiLEERc/bDFHaz5GSJvizT9OXNQRJLrw6n/XG6Iv5f540rlvqp1ByB
HvqS4wVzP5Rf9faBVo5rdE7PjM/ihyxc5SuJpipACFALczIs92rdPZVh2mlNCgR+
8QPLM2SVFAQMEsaknuD10vQBUPlk2WtLEDIktc8Rjoz5oijwCGfRwIgzXPviqCoe
hk0GBHAtqsgkaUirI1U4y9Hmkk/2cbJptHlZ+xYuWuDovAA6/qw+PE5ou+PjWMIP
UAaDqM6R2z/mHmJy4er+97JK8/1mMCXL6gi9n3hsuZNCR+hffstenkuIzRZNePLR
NxD8Z7YdVHdd4i+kGuMZlpoeUA1EnfrZOReL8YlbdCuhZSAoUXB81qZ5yFhu0kH8
IIYPvUriKSGFnNxzvtCmLE41M091ay8jnXUexfZbBPLFq3/MBHTdv12s+eG6pv4o
fvUwAER62R419uTBIv9AdIXuUgZlF3+Q2CDUMt3wQ4A0dyUN6j+76abZ8WbHwv7V
DJ6tRxmsLTQ1RAYO611ImDrwlnl6a3EY9qOIUiBhzOe+DDddwd+f53D3QmxTmQR9
RPkHnp6RdwH14ldETREAwX4x9w2gZs460WBZ5KPGX4iMS5Jo2PGPT3YshW9fZ22L
lQUuNkEL/oHutSQfhLZnkEAddkK5UROpEedYlUK/rp1wbCguUyjGMDitxQ1KqWAi
h0G/mEyYNOWlIDLGLF2ffR/6DMBJ5cuEsfPX1+37zgZuuGA8zFLa+uA1RXBEPrHU
o3PaCGR4Z6jKz1DRBm62FVO27UIOmjwONycYfj82iz5MgRjA9ZkxS1V/iEB7i1Kv
2LKMIwjK+ZpHKBELnzUdgm0xuXJadY0Ctlg/S+0CWusZl1zOzge0bmn7GCJMQpRy
u72nWkIAl5TOyzx/oPzeZvcw3s7MhHCsNUberHsgQxPXyskAfinOvDbxTJ+IDD9u
wuw16Rbe93JSgMFUCLOsbrOZiEglv3XnX/luNDSiLruxN3cpRYQ7BTbUnWqPRO5s
ExxR0uX4Y2I3pVCYcOBEa8cy6j96oVto5g4j77pLdxUFYYylpZQGflixH8AYSUkQ
EPmD9NFwp15HakK/yvY3keVWBO7o0ZZKGC66RJlCHoHPkmSt7OvaHRFOEuMd09uN
i4hF9YeA5iOcpphQC07orc669kholg8ANQLOx5I7YbQ0hiqn4rhliAznhWQWcVM0
6nCUoNVZv1fYeFKsxKZn9J4/x+RM0SRO7VTgOxBHW5HE9zX3pxy9GJok51KPwYNu
k7g8Oub0wyXnx3cJAOfsHkjCM7D0tOas05ECpjOM2DheJY9AK0vbZUJ6/Eu6vZ2a
n1eNjDS5xUgbGnIYGRWtwQ45AuHAhpY+wWfWHwDmED71S20CfRuy1USADxO2Fh5e
A0HqnD6Pf2S+77EcX07BT1iY4C2u/fRpn3EovJ5lpvXuA91LSPAMJxUFjpVFurcC
t4LVbjrx6zcCZql+Cq1Qt7pmaFspToW296//efUHgSx0XQbSICFTYNk9YALYuohc
0N1JwhhgSu7zH4sLbwpSukZ0wED+Tz26P0HnC26dR8aQiilJ+L4qF2DFmTvYnFwN
dwbzn4u4nUfSR3mJrkzxiDtUD6PXscoq8rPs2uK6vHQrIr1k7Ga0qEtPgkWtasKn
gkip0y3adC0S1p6p9iW6ZMYYItiNhDPqcM2tJd9PoLeMOgNHIjjFSWnypM0PfZxb
0fsfFtKQwtA+skHQIw9B6KcZwqn4NsYJgOy4Ys5w4tuzwFntou/vow8+ZvnL8ynw
WQlFmR0TSt8w9APN72XI+NRPM+7wV5q08n8cebal8lXq2v2SIu0jgsezkZukiqdo
DOphfNTfyXYgfgjg1qWyP10FZa+0zLlSU9tGZ4mwCRiYphr/0Bi3kgIPQUO7ci1F
RUIVoP9ozBwFIIUiCIA8y736rYIvLgb0Ch3RAeV8yIuxde3L4JNGpimEGgPnFRy3
A5syeIuipy3yx2crE9kcZF4Utw4kP3aAI6cKYcDA2TJ6FwEBfx82fO3j/d3KCbvK
lXM9zXdPDJ3p1a8udsXiYjH4CQFXxj00AWfbvl0mZd5+v04AvgI4eRXzsa9ioI6y
AJVRVYcDcgWwXST5+mF/5/QCcit3kJt1BVvZ/ri0wvmWVqHnJUU4wWsFmAuJDWqO
w8JIIunvyWsbSba/VtcAuiQjn2bWTx+QBdjCc8geUQkJqZp3z0+JeXYsGtZk5MEG
PAnAc53z5euMcvkE0nYH8nnBz+A7TJKMMsfbO1qxp2fIayh5gi4lXiJg1rs/2z89
+XOO36w/k2+CL1TQc4hHTkSCwEBIKo9S/ZaxQY3NeXkGH6jBlqijM5DakZNTiJDr
R5IOhqBd3sOBP/dZHrp96u0QGSeuUt8Xwm+MLkjfz/6woLh9i11AiteEqn3ShJGR
Q1INEz2UegSU94jpJv8raxpGBGa8BBvbwyTw0hiT/h4eek2J1297tKJOXGtQcRfQ
b+cujW7+CF/m1FXd5Be0TtYUlKT7uMBSKeEkCYOp1a4SuHdvAOU+yeAHQssI5oGJ
LkD6Csw6kA8FocnF1AJ1MrqtaYFTxST3kmdrlD8Z/ayzutQ/1DkHzyFXq9LvIcV9
IR9+e/qvqvt6j9jKF0W2o7WXCJ8vU4rXsIf+aJiF3zeVTy2Q/+dl9fsPs7wPhVNK
EquxnxmjVLLQSJfyTLyFjt2L3d0BJCi0hIx7H5f75I+43jhHceriMEmLU+4X2h16
UH7BTm1nnvMjV13GCjKl3vWV2bsl6AvwRudi6S64QrspToIADdntzezour077msG
r4qzd78N3mwUHqT30uPihlFNPH1AvqTWhUWZGj95qkWL2wisqJQqPa+HtJrk95lL
Rpp5oHNpPIkYm5w98tf6INJ3cnoaiQ+BaBDSa5X/8z5S4ynaB+FANKtBomW7GdKI
An7i5EcMgQcZf8o8qKZ9cXoXSdTGvO3gvX0x2y+nZ9ESCpC6QwwRf6AifnRJ+jA1
LUZm4rQrgUni0nZmO4Zo+EvuhLWhUYganjE9cWhdOHX90DL8XNKmjI72LwsvXKXn
c8ZQxH9lRI/Q5ez9UVO4WP3fmonJ46p1gFySN2QCWwijZP0mPett+/vnPZ98bqw0
o1OamiQYpQBtQ65hUf/V+506Ifn904rp9kI17xC6LtNYJPIBig1DaQIQROl2g76E
QDzxjunlCgZCXMDMBR/U/YSiFfDiWQ7AAXxFPNM12alo8rnAanvkGr1+BPIDPh9F
vPLz9L54XPYuEAwtgPrHmBj7gyhv9JINGbvW1yLneQrHVvLlxq/9Es6j3ZjGdzD1
YWfSItSQVDfQ2sJXIefJHRwJoTXRRAMJ72IxYwFipgHGJN+RoiW7pi3XJ8Lvn3bO
U9zBBYbIcQVgM+N04aGkkHBj2mM7HJxv7vUApIdiNAu8fl45SZd0cXRvH5x638aR
iGVeetoeEwbr/1dVHIuTg4olAk2H0mN921PB+O5vaXu+Xpmtivmi1cyMg68vQGCj
tXRBDx6cPLZb0UK3g+I98LxVe+hSb51zjwFE1Sj3WvgL5kOgIxzuuKRv0R6TB+Op
lRQpcS9iHTqRTldaBW+pNdCUuGiWgpmXZBusnMNydsIYzpUXj3X8CmRfQHlmQAVd
LLd3KuF/ysFqsmWRKinzHK0CECy9f59O2og4mhUkxtzpdhnHOGcYPmBwtuznwJEl
OZTuCdwnq0/8m+peWtixKjA3DxMMNMNxNBUJTztCk0u0+zdOiaVRBTJYlTuCUvvm
5wv/J8RmAhcRBhZP9FUR621++X0NOfzMrKo7vxpeZmITJh2iVhNVBNbihu4mVosb
mWXZ1HQCHRCUrMQozPOlSIF3P3Zj6pifnWNlOvzjLXiTG3ILnkJfduN8N50MbQ8g
QKz/d4lorllf8FfXRDgePtN8f1vlMhIn92naBvwyUr/3MnwoKkw1TESuZyGoRO1h
pCXlQzGPTJkVVuPefsKkmp3af3F3ajgNaAvZC0H9ZMZxfBSz7rnInadUjIqFsq14
VdcJlcSjioGKarLdeKt6r8Asb1Wd2fkdTFMPUE2WUqXj+Gk2IQnwCXJPvo2I7Ztu
mW40ZNLZCEjd3J+iA3oM4OPJ65VTDNfOUkaozsW8aPxpHp1GM4+b+OUCEmSzEeml
oUr+4L8UDqhFUbco6RHwmX3EwfhlZYfgAq2NxdkSiMs81oBh1VAlwqMDNDPige8n
wgW1dJTqRnEV6Dhpu/eL+Kt1mP2etL9nqzVzasr7GXtcFx0adZpNtgLo2T+g0uJg
1xZx7hc902tclOoaHnVWHs3WZCR6KAV2YzlO/h/yVtgYrc9pK4lUGlGiIfQVchyp
Dap6nEVnmRhk54WeV8ij+KWNURDDibKWn1i9t28z6SQ95+VYzIpZ9IKiV1rxyB6r
hOl73rT+J1xeflLYmapBUwHMFRaoR2ZgviOIvvoNYU3U50++WKDwgoizaNV5iWrz
lVsbCxJVMDZHILGa4z2oAES4b6TwHH0ssKOXwGwAal46iiWeolfPaCILqYogduwx
lvDHXIsbzfXSobilFShToSZkCQTsUd6EyxU+oJNjK1eCDag/kF+HqpXeFYXKB3Ze
o0I2JkvtkWhKNw277nI4IBjIRVHi+WDLFPCmG3JlF9pqZQZfPbrnLidmTm6W+jfg
K3/b0OhUunBkvMIfL012W1whrSy6uu2TAje3dnTWjW5WsPEnbmcHazuFbVb+r4ON
4uPnIzL5fS43Yp55P6FnAVB+DqB8entioEboAAEgaADNjhC+l7pWCDLN0QB4p+Ms
vgj1oBEA9Dg53yUOVr1wJo4d0O78Yv3hZTEgheHUqNguOG8dYWvMoOgqKw03riyJ
sC4egTmbF/GXEcbyu/Z/+C9z5v4s4iIS1O+U2qVtEnhFQpUd0qiSXrTAj8fyUtEo
i9gSOuGvH4bZdUld0ppse1TjEg4YMwG9xqAVL9QCsFeAUxqhdUPh43ZsmrbtmF9m
80SFqS0unOmeqvzEXisvb8pKLkCGMztNis6pJCCchSnl0x/PAUfYAhxqWeU7VFCD
lMBmegfuPCEekOf1e5tH+ZROzBOfwWBrd35OF1S3zoNw1ocHMcWbdWwG5Fok55ns
qadYAZida6GxTCc2HVa+3vGrvHJjEcGgH6RoKX8YcJq1xghgXuFkH8UEd6PlrOKQ
1pVBGragFBHcfvUnCVYX33jt2BaUeoGoLUfAkBV9GyEjeTl+5a5HSt6ExykddK5F
a4hrwdPLX0jbrbvePzZybOSosaHYWaqUDuFjIx4IlfeQ4aPYdLu2rdBDS8NyRhG6
Y2WzhZXI9Kr2J6TTYLffK69Y7Ix+RVjoB+rPaPVCJ/yuEgJEfknyZYXakTi+SxXQ
uIxWh1cmfDomSPCOga3eZ2sdWdlk2BZd4SdE5Lo87jt/m0QIFipZy/o+rTTbDSwh
XWnWuJC+CSXjzYAc/sUhpPo56H1mD0tv3CyCWKBD9Ku9IaR0k+fL63q1OZPzgelK
Zh4yy3z5U1dwCe/5IO+T+qceEI7JZQp3uQlTeNqGqh5L7TrlMjZxhUYKhZ/PSETC
i/JKTT6oW8h0yXRtrjcaIMS18VjTcLlhDII1zQrKRJLOQaLz0VyKVnudKd5I1IFO
engRODMg9pb1iQ2R5Mhq1SNGDrA+AEckI9sGhMWySLX9nuvDGGGqa4OARU4jR3KA
VAUHaOXut8sVRpmMba4UtXeutr+Pq1BkQt297yfHA/8EPS5PSBY/QbDd5yslAnTF
tsn46NVHh9SEcG9mrlxoXHAc3sT9d/wZVQh5c2iAsOzr0fo9nTa6MVXchd1f3+W2
ihXu+cdECWtdkxQ0Ug0BTEk8CD+azMwmHocCvfHcIgYbRwcfgMQgYdAGEOBMiYkl
xpBtETWjtPSOCiMNxlECJlKa7GNGQfAJ2Nh7wbjivd2SSufuY+YBUinK6RP+/hPp
qPeJB7wc/wmlQHMH6hj+j+0LO67AnbFANrrui6AYC8ETyP5r51a0wPlniIkLtjpO
JQ5z76NuJo8UccYNtrQ0ZI+qSvJ3FqdGvp0yEwIwx+jyLouPuA7o2Pdi8fBV2DIh
I+bPaU2h70cF4sDVki/YjStnzRFfvnzdXomUc5nR34ryibdD3b83F2QwZSyadWCb
WZjDGp5RYb0QzQXHsl5/m/MT7dH/PhZbWsvfKqClH3OBH6J/WTO2ohDmo+R45vr7
VoNqdbEYhaCV9UuoRleBlaL6peVGFjAm9rY1Z4mVB6A+hxfLCPAcP51EHr3igw0P
yG3/zWlohUbAS58tMcF6LQCFrh2KWCAlLln0+K43yZP+bWAz03La+iSJ7SmgZfh8
ho9ui1GWQIxZYTTBEClikFSRj5rcYZWVg6QzfW3LeLNZwEYeXGJ0N8W4Ss59iiKS
rqjHmsvCPmCyjElfaTS1kTLurab1/z5uM3xJyPX2HxC//g4a0I42QA7u/Q+wfX/S
9/ST6rz9IKIunV5YxG+DhmcdzNegjFJ4fPdChJqBy9xkg8Fwd35oRr+hQBI4Ys0S
YzBvPQO5OjCkibGHrTG4FdZFOMqe5B4ZCTuwiq8dF2H0UhPWOftkUNrU9ann7CMq
Ds8FnARUJFWPMcAOGdzI+b+eWbvfoy+lTmFPmBVjoiddqLUJxJCbdEcR0gFJ3zu2
w7q4duVqAXMC9wMHG53mKNWS40fySXW92Y5O0BVAmFaxL2WQZenL/PV92JMaKYre
6GpWSXS83g4Z9k9z66MMNzKkn3tJOLs/sPzki81ClVgHZh/B0wrzeoSZYnzx+jxO
GWjDPoR3HCc9eNTHQ65miIbzbzWPYwSNsOlb1B1i3KjYPs4LJI770W8oWSAz1rYE
VeZ/SmuQ0JwPvw7YXAZsLt6E4EHSdorw1B+Sv9V0jTCCb1duMEIbBGYbGAmWzZJH
vCDF8QnUPazDuh5KfUH1YlfBi1e59EefJiK+RKk5w6tMcOPirXPdSs05DE5wc4zz
RbaMs0Flxa8+3TI5bBkpEmZ0xxEZ2NN3VzSqjhqpW3WFu3hzuTI0AkmbfRfTYSA1
f/d8mZ0Dxi+hFhnX4FX8ft11iO2kMbbaeQV82oGvifMszCw9yeervcOuQ22R/k9x
Rc8Md9sz/gifg2V+UE+kBdwv6ai9S67BT1nT82Z7YPtv9dNBFFMrFHS4macTRa35
70Pax/4g4YRRGFwR2hbXGYfC0Zc6bCNH/7nt+o8j9GW2wb+sCgMRR6vbaRWd0FXD
vq/jnhkjHn7Qbtf8yzzXSEQDlFKa3jZS40ODRzE5Pgg/Ynw5wU2mRuEg7hoDPSMK
mcnnX6wj9JB04regjleX0OXIp0A+z4iJ1ALc6knw2ZdAZ+TCcIfrW3EnzTmg71wc
6bjcU2mhPel8kIuS1pYhp73rpZ+bgegGEfIPI/Vr1V1T047JwhuWsPC5r7YTi5vG
m567mM4qP0ZU6ZF83v10HUhme2t953VV4pz0d0qd/H5PjWfDUUMzWs5EtFbDn4tZ
0TQrvlumVh4fBCPpPnVjVpASdTSFrEsCWUJeu/G90HBrnzjIob/LODk1awTnlN5b
Q0jwOjtUEolM1aWkZIhhYMQqVgh0n/AZLv9P6hoAksn4+MB79r6CZPp2biJAHLnN
PALPC3K1fbtDN+R02x1laQbD3+FPI/3nW2eHWOxBwrp+NBLOu7iwz5WglXISlMy2
KVl1wBcln/JYXdaIym8vKf2Ue178QtVAGuXe8HYZln6dnRJh4/i3wKdWMWpsSfsL
FTkgyGe5AMIEKC5mLqAZts1Vn/SRe63QrOw7b3YRS5SO9T2DWqa73s2a+QChE1yW
CE4PfAbgqdqk0UKICQ7PKpjKCFBWL5bUyH/de5pIUoXZOuSwk3smr3Aoy9N4MqMq
KcsAlKcZR2q6XvZehtW739Fj1r5E5nswPQmY4MvYQFBf9hRrE747NAtfWQRZ4xGy
Yj9Pi6EJJwazF4Z7Yms2fv5eaYWK0SiJcYxZjTtUXsARvlG4HFMWwysPRtsj1I0b
80Ft1GXBbmHrIPVImbUOhlB0cR/db8ASPmuQNKCiiHruC7yg8t1QM/ndctGatxXO
+8Bz6TBPd/4n9H4r/BYlgkI0h43iXonFza17Kk7uCD+aKB3fzeX9Dp6sxHgbfrvP
QpdS4X/QrgmLZoWhaMiP0IkRNzGv9rMTszWAcjFX6c7znFJ/qE9lBHtdYP+DF9Mx
MjSJhVIhSkT8qaP742NHgisDlBxhHyCrst30GkDLqHKB6wSpyPSHXCZHybcsyYoJ
b3OgOWF++Ow7JCaIYrsSvP7jtL+8ocsaL8H3Re3CPU/BBzcNnRHxyBGYsr2tdlXx
hPSMYhrANow7ExZwaMj1y8WLlFaNGHEeXlLrnvJnV5YnbDxQQXKD0HomM5iW7cag
stQC7oFtiqS3HT4sG0zVmw9Lrz8lB5WQUu8HjFzMBURzBAQSTRRIXtFsTTaM99Uz
bPiZyM+fbNH/p5MoI03pS5QQ+mZImrgm98WrsnCRhJChBmxKvrgsKPlElJKGkkT8
AL37kW+vF1YVqryLN5v4xjvgTwp9CE6sbodHuTem+HyrBdA8vecO8uvkyGG6sNUg
OClkXDVjImD1IqQyfUu5CHyF6FlMblDyJN9eGtHz2GC1cAIqX2cGqQ5XDukdK6C6
td7XR8dx4vgpjMBUJrCMyhGn66G+ZaP9aXTLnz8mjwl3eWdcqPcePJqnQM+ZdlGT
TCsbKUOnItzI8PWQx1pBPa8GUNC5HVKiz0LD/BbePMLjogfR7zuVWldmiWYvSNp9
3jg1UCVQf+LerJ+gbdpP4yHrz2Xm/WtJsNrXjuG8x98BqY94HxefWHN+q305qqHK
es5Xq/11X9JHXVUvzOpVv+4C7Zoo7TOvq/COCuqXnunwX2fSvcmInK/7Bu/gVvP3
UPr5oom/VX5JqrGFWgBiw1O36DNVu5aUoiwjQLlZUy+N2W02TXysmtubWwuPk3ln
wjGQlMynyYfRxCTdmvzOTSlQ29Vl7YydPyIaAZoCkERQ3rPFcJgrgvY+52S1gHDe
8Jf8snhongd3a8xzYW/T3Bdc91ZG4bcJ4pFCA32CLxq3DvKw5IwMazmv8j2HKT3K
fJDY0lRaaW1rcJlj4ITtvz5VmnJarCI5RDKA3G7DwAGqyzpROaPxTcMx/vYQf6k9
JJyzHDtbaD66DDEEfKgadbxQEF6R+ekJV8s/IhkBW1Hfo475+xQOiS7kiwlbry/z
jaB6KaUz5b+Z5yuAmOE1hGByIrAOOe4/8CS+wd1ZrPm0Xu8NFVe6JxKLwwVYduxI
HXGmyG/0XssvqKVEDAYu7qgcU0dF4zVbGxuhG0u2k+3AiqmixcMesswlS7TH0DJM
5GrJ6f4v8Js5Vv8TGnPMGOlHEAJI2rUF0O9hx4NOKMDWOe/9VWhAMyMZ0+ojsnAO
tMjpnRBKJUoqneaK7y+J++86XhsU5xlww/n7INfgCRjh/nRurdKitgm9O+Sh4uNG
tw/9ePJOoO+vCqnpF8FSl9+eL/u39Oc2JiqSS8uhu7EVx/HEHgzRfx/HZmIsham0
FzqBiq0uc51cHYXW5+gIqBU2TanNqCh1ys587qsPuDachRaCZqq1IoXnLNbWyDFY
38Bj81CQbKGsu9XOIkC8whRibKoWeRjpfJXIHLP44jz+3ZZvdX5Hi2PTnoFGulyZ
kcLWbCr4gYM/7KkGr6FLEA+Ny3gSfIz50BFoWMKRRG9RUWhb8eR4nU9UP+PJuaRZ
gZ3YaoASmkjg65GWe7H9rQ8OCsu5GiaSfcEPWyw2f45GCbYUPhWpejx1TQfEMM8Q
u/ou2d8ilZotBeYje+8b61KIus20DZEyeONqiOVJlfEZZj3x7NDr5Xl4fWU+9aX5
PYMKWyTDxtlU5P1ZFaKy6eaUCDGaA8k34Bw14ZXzmRmRo7z7kFh2hkAKbIsqmwoo
5OnlCQRgdWLkceJ1oFMc9YzXJxFpzQHvtZi/QTQdTRWGcqSKKyJJw67EDdnTdFaH
AswOeZKANDYoUS+YRO5v1tXcvNPVkdH5bLiJ7RFNEP1M0jTKJ06V4shYc3fjPoNY
Henc2I1fhV/DpLIXCSr5NsDRLrf4XOmts/qUihFbkuY0BaEbTuLXT4kIvhEPNTtc
sxOWDsx6FjWgxLgfBAdocDrNpUZFL95jMW8FhIfWly95yQLAgZcG1+Yfk07jNcnG
OBQr980U47l81RMcmp6rBNi3FJ6+yNLSVPeFWGPESukOiEMzCJrxkdA53RYTawhl
wLwJvMmDYWXbbshTX+MgATHKWC0/BL9PUD9YCFe/DYmwAhNuHmRmMxGX8F/qUaOG
H4Bj+it164zfe1Mmph+Z/6/BVZec+wL06fedDx94QoDii5WyiHIkbiWHN0z55iWH
eo1I3Ejv6W9ZpfCC1a+ovGEtN1vpdjkzGqz9ZdY1jhB/0zsd2zIbNab3LYRWkP9R
Q1WC/S5jpuowYXB/eh08EjZ75CTPbpUbozUthRTA0Od/dlqYuqnJ+/nbGL/GmSig
jOvcKih+EI1fAWo1e05KtgM0KAsOy1i8Vgc9liaccPVrN0UbokG9UP14vR8sqrRw
UKr6XziZxNuoIxv2iVRMHIgMqNaaKvRqe8uq3MrRb5ekzH+HllGmIY8IpLmuzFgG
7FjHh5U3+h5cjuY/k3Ie1FHhYBV+8/Ye3EA9sxheSwZyXKrvREMbwKCNO3oo7pQI
tRQSwsa7WbeIC+ZtxR7OneC+0INu237CNt1Fr1g+m5tsaEl6JvfRjegAFvOJFprp
ghcpwQ0j7zs4RBfFMVUdJ0O7yYYxvWci8HJiFccNUMZ0G0UWuzGcPJUbBZ8JKbwU
iHtmdqDX4qaZEiaVCeIdF79+j+AASsAwn3y5xi7IbFfyvES7E8WAetVhA424lvYo
pTiek/FCIskXVSfWC2CHvEKMKzGKu4nIP3N+A1XH2+UJLJbluR3XovaqyywmcsPA
Eg99Z3YYhIjmrE4XU7cGYGfp3fkoV2E1to7cMfojBvcwac8YkeimPlBUTMt6FKOm
2S0Zw+xtUMKONl0UUmyQQzwFaI7KFr9lDix775fxS21IApzMCdsmWX+TP0LPa3DC
j/QrdW0G0id2HZgKekyr6eQF0NzchVI2WP0EwT/PUcJw0zTjKYSYVTbM6YHIwuhW
sSYRQxzpIGA+JLSWc5UpiwRn3cV4Ig/Vep2M3NBScpXDfPcS9UDFjyngSxrrz0mH
w9HsjLGB9OFiG4jG3gPAMkYaasuPB1A96oz0NrUmv/rkaCfrfqyblnL3B2owQ2jD
nJRSW6pJs03qMLF+I93vjtdXPTTpt99t78kM8J/AJShBgzYDd8OJY21CZhnMNwms
G7P1gipgCS1X0j83mVpcVbsNnxOXcKjruy35AWZUC2jtiYHsULQwKST26VXRbrUq
ZrIkJDJ/gtexeFKaaf4rdkQoqzYqkkkbZ++4qrSlhQluVR8UB+BcyxhnWdTBD5Ic
pK50PSHa2Tj15O+NZa98TP6uE6Rkioq/vaEaaE2znDZhGpJjwDrmIwLk5E21hj6+
PFiZ5bAVBxo7fjoAF/+5l5YkZyzb67lUP9jpENrUGF8i3kgMJQOxWozGZG2wU8X1
HM4rxAsbro8mMcKPhKlH2otFnOb8PFlS9qf5H62ssECSqZlaZXIuje8OXkWGe043
9Rbq21MXLFxCT6nx140UvhfyCsq4BFWjthmlYWFVJ+tCNNZyt8QoHBOw+7pzAkZO
/TQWPX7D7Ooa2IGWylgc7qzUhLXmyOq7p1XFyF2AqMz2c+abcDpNx9Y8XDTIdkXF
J799jxtfDlt82eGbxh22y962DdoBJm1u//gDkpUt/D3Kwr8JWagaSqWZM+l/KrAm
06YD/8UR+8hh1Hm87Mv3/SuDpi9Edx7zDlbcR3QJYbpdQGRpEJAxpIgyIadhpzAW
uE39d3nxBGNR6hqN+FkbVdkjVkfcQe6jZTwjEaWRUaHP96c6679P6wZ9y79ipdUy
PLDSIOBoCC+Vem/JsJM8kDnBfFpESxogOq6OKPcr8mxHIoN/y5vD6Hg5tDAovTGA
/zil7r0qmUVsSPF8nvnD8bnNgPv8qsqQnUcy2anROBUWRO+1SL8s5u8yG8pJJKIR
e7hO1le+boY5R3zGBqjU19GzHt7x+U91WGUpr+jPLpZ3TaYR6lSbYw0tvRVsgg4C
QNOlfcB/h2qwe/P0P+FE0MaZOg/QhiMXqtKQLx7y8XdxyZ3JzFNcs15xayReHN3h
40haljyiAsOlsgVXRiueKzHw1Oe0Dyn1/nCiaxNbPQerG9JDFiZ4/fyRAWnZ7rOz
Ij/9BNlJPY3soAuc9qUfhYHu6lKwkaNlerXwqT8oxn6AG99AHO/Fee8lPm8Fowex
Jti6slmvOg4ouEIsuWXhZEtcu+qbEQGHcmgrYWV0eV2NPUoG0OBZq4snRlwocfzO
jNEX33pup/086nmhfuPLju77/B/VJJ4ZRLPGEidvfTc4EZfxX/9pBHWaHeGbURI0
dlOMTl9QcCWUrzgC33butCJ7fGHKW6+Dcsh8FJdYsjGMsnPV1IIydHrSSz9ujjiq
wQgpWLTIwRGx3N/MgXwACzNK0KkyH5ghTfrBuad79zAdWWWmUXt5awD1PY92a+WJ
NBqV0+ldeb2zfMrg30cKNJz8X8oTaNW+/p/TamF7q9QTALN1EQPKYO2hTnjqNJrG
ryeMQ2sSGmsMC4LjflQCV4vsqLKx8sx5qBRKRwalQxsNLOX83GEtLDbCfFj0hyiQ
FETWJkaTRCTXGjYP3yTRZGeZEanuS7d3wwKwpI5UxElA1UJUZCq0D3ziKINDtWgD
5ggLyTP1Z3nrSzDEfVg7BrKLbi2QxRqAchJq81EmpDRUcE1RKXmGkH1/C3lE7gOx
kKONB//PcFqd/vVZjx+b1vAY6YwcxY1a1hN3ECsPY5+uhWJQKcRP3M74ByJ6SC6r
H7EsGYS5+Ev5GikgFt+00VP10JFqms+opjFVYYQvnayMAu6Eh/Lepls/+VaRdpTE
WDeyp9TRoOWoMwZcl33MFcWuZnuNSm+FcWcUBvRFgBxB5gHuyjH76kh3MMPt3mvI
AkfG9ZondO5jrD5GMqZmfs5/mcgQbmIXHSju/axC2Ay+jeaY4ct+PCq3xqH1vP5I
d4oN6cHkHRbBRRWLbB/JdfSNg1vKEHoMEczxyjuz2q+TvYj/wc/WY8GNcgC66nzZ
HhiAi32iz2HQE4fZ7wCAMc/MK6faLWrZahRPljnIYVnF7/KDb2dcRpiI5+SzermC
6fPh3ZM254G8l8zg1vS94nJUOfD9WiKbH/pEO+8BXbxaMgEDo7d6QauEzq8qrHJM
2bpBrPrO24IPXW5T7m+ejJHD8rJEyNtOeUElXqrv2/IieyopuIw2kPcgRHxMFNop
tD2W3g/Uy8z1S14AlFtzC/FEZZocQf9t8vLR3TfZ3xtkQNqO0F8Mf9xooO4SxyoW
ItT2BNGD9SKqbWRLO50dICybA4Gfsa42SLU+DIj2YcdPJlBkvnDScDOzY/oxKWOe
Bul57pHZ44wDkdGhq1iWcfLBsOHEqtq2kZDmhj8R3n9uo5k037nZSh5VJYYr6eR5
OM3sL3P0sZAzfiNew/pKByXCl6+tq1vfMQ73TM0bDET3oR5fvLQlCBqpvaj8KEov
ZZc0GDEFWBmI1/60y3SRIs9xY7HF3AUMvMZQx1VT0zSgzpDmwEAes0L8q2Hos1fP
/hSCM5LgyBBqPqbKMWj3SiEAIdtG3y9T37bUIoAM5zWp3GzolhZbdFxN1zkheg2r
orFq2p20cQLP45qT4SoGo3mVF4JivH9NMq0JamhqJ43sFJ4wK9t00bVEuLNE+z3m
Ux+e6rb3nEQlXqjIbArHG3CRE8V43hpg11znYpeyjNGCRru4HpVuh9M55PVyV05+
EfGcRwBDz3bLzukpvN0d80L4DGX47+itnvANmwU4NvDCN/TQijT+mcrkn8kbZtVq
WqU3r/dR0oATeT8n7kOiamdKZLC+oCTS5qsDHWz8FQMYm60m8/PZc8pSgqeHZhVd
IOxECnUH2QERSyTrwQIDVxnRkPbhE26r7/e+acsJ2E8FIBz62J8NzePn/OyCmvEM
rUs9Lz0uPuzH2K4QhbGrl6/JetJ3ib5G4lY0q8mzxDoYb8Z+tYyN128ldRB7DdHq
lfoCRW1glyFT4Aj4B0EZf8ZLj4UxuXsmroiSt3jge3hZbd/Ap8ACjYSYj5sx8bMM
u9cRFm3PhTEXHFYmnMlyjAUIWDZ6MHOZ5CJskIc8UhCVcjPwLZK6rNdfAvcCqxcK
fcogNmykH0xu3R7iFPGkkWARwSbBBQeiXiHv8NClzTykZ7oacxDyT4xuZsXnYF4y
p1Bg4cZrTZHsPp7N4fHkHBrk8FjDN24GPsVgxxzPJB9ocXovzIjMvd3KqkhTnLQv
fxoddvpBAwxUOvc6TTJQfaHMjUsYMsxLwLFUSFsxYEqrCkA8XvfS/1/zvlLZfo5d
+RzEzvnwpnrFDXGRsJ53hS3QZJa4u2r72KsJaAYQ+Pqp4pXoXAxlLmNTlSiFB+Ku
rfodLzZYK51eQCpbZoRTtTUagiZBGXSZ9eLUMdYzGT67BRlqCLqd0G4cM9wHc3gs
QS6koEJw3ARk7vP12JIKer/e1jdztskJ7sbWShQikWOpqCcfbqGM1/8s2oUPgKca
lOxv1CGtPdi1OZIu6t/6NNr4lSe09rVzIrvYLmAdcHhOCw6S4mchw854lYEnJG59
9uOThtL/6JnrCrehWHyKasOgCVuG2ww/1Tv0iTHisCcp51qrqcV7pbuoxRYdgo7K
iajxPWgGxP9vngEGsNZZBchNX8puv8oMhoeJuDZaHHUF5MeuDiCXlviDouEk2ILh
F+fBimDw3b6TE2Ghu0qf85ftfZYdEbYJ5tZNfT9+H2JFlqiE78QdBBQmHS7HHn7V
TFpz4CUwJ6EYd/CsOa3SlyIT6WVdHfIGvsCHXNPj4bMr4xVBui+Oyfq7BSqjrvkl
34RoZuXYJDmhFLYF4+lyRcMVAMVWLjc+d+a8EPbI5/LyNotf1hnyf6OclToyFSfi
PPL1jp/5ZIeGjLwlsVMoj/UbYyJ7qZoP9TOXnMKASvv0srihRSLvOBobbLCY5Evb
/EPYzcBGLpwgCCKwP9vdGC1JAwGvy+BS2UWlkM2pX78r+dBnMPbJW+S2lBh0DcIP
KR6mBTs4VQJoXhSx+liCi5F/utCbf4ZL62vnbCfIZ8v6L1XH2GjVPtwuLFOeztsv
5Qz9k0CD+0peZT5TBEIwlDEbkISZ1MP+lbDEQyMx/8fprafbjszdFSGnvlYWgYh8
eaLk0ZcC7+fznq0pSMzO9+lsq+sbsDlpMJK1MYKaqmLnoxIw3qIc0HAWDIHl7JEs
sUeY/ICaX6HpjNimnr7goHrPflzQrCkAbH4FmXYxBspV7vtQqQBnSJ63WZ/q0OLf
MaEHAeWvu+dlMSINKYI2k39klMeZrXslICwovz8qP31eYAGywDV1WtjlK3VTvcJG
uD2goJRLW8QNQAWfBFpRgzIqyenHA/zQnh4reofRUZi0TOwm04MWlE1J0wYmlJca
sz9Nk4aPjo4Ut0JADAsSVLmtnWksN0CLRvW28PXdXeI9EcKNcBtLneI7ZY2o0U1P
9f/JlBKIW/TlSszt7GC2cTqIcq4pgfY8BOZpyk0GCXNarvQMoQLG9iWqizfM+5tJ
7d7AXY4Tnqyj/hQ57Sb+SQqnkTbvjDW9FFwmgFVCh12ItQ21XW0ozRm4dolCjSu5
H2pnhiBFIL7XCiit7mWQqeOODhphJqzR9j0IoGluO12kwbwtBoXbsCZ+lyyKLkv/
gcin+gGg1OCV5IGaNKXfgyHFDtFGOjImERSTZYqA7mA8LWWpbYleSZit0eGgbRWl
g7CBtmDTbkCnqtdvzgUJTh4d9roLedRRDkujF5UDz5dHQYOhTTQH6OFXXhOzmBCP
BhE7JappgD7KelcXSpRvuTV/p7R0uI5f6OczNYY+5jShboMvUI7jEJmEN4eZl8nU
+3WMSAkJn1+ED9UQqbQaVUB37rJrq8Nw1cSMLjZCTO8+3xFCrbfdER1GJrZoF0PN
yM0JuN+HnE0qOpAFTuMgd03heamtPC9xpk3y+S3RGRQqT1HivJBqG7gLq4NvBU+2
t3ItE8zj4nf8K5tDY1rUWfryYBDYCqixj4iX94Jgi066TjvLNFOQ7UfyC/m+4j0I
/4pbDvujN0VC+WfZCf4Lf/CsJEf//9c34ALLy7/s61n/fIPkKY5FHJSmWVKfBsSw
OwxhVxuqBnU4Q92ISkSXlfGpe8PhISBFSZjVSA6g+H8U/kdNDIEzxPGVUo5C3aoo
F3lGizKYu8Sju1EiX224t1VeEgTqdPDVulFW/EUUmn8ppwW6PvhqHuCEH9SXmg/E
C7hNl7j3zi+f7jdSMVJMS8WkjPQ5zPmSRqZaOzZQXJaZB2Rm6up6DoL2No529qW+
qYxxKOPOn08rjLIA1Pn97OVTsA4Gh2E/ZG78eaCsZP9r4clw7LcYgNhNbW058w/X
8TyFTA0lpxT93axq2GyYig+KhY2M+LFaCeswNJdCy03/Wga+TcDLFrt+FYxBmOFg
KTWT15NovbdlNjaB4UG6i3QZvMM1/kaHHF4etJcvhd25/kt0lRyhXlJuMmgoSLtk
ZGgeJjUTh0HHi9Yl3KwK31rUIw2CTgRIX1955IUa8gMnJe4c1V7gfJMmMc9DpOm5
zm+YzZoTArhgLSvt9hpppwvllUPxCHm+14sBDie9rfp/KPzBwranFTYD1Sf3Y3G5
NV/q5j97+WuXa7m6h6WEoXsPCC4lHaG3oLF50XHPfgKSi93JMjX0F2QQFM7bh/32
0z8O1lLiIlus4z/wOWwij0iThZtXPXNLXOKh+KjOhdLv16bygBUGcihcnxYVYwus
2yBa5owEsIVmRmnveMXEsukmX7jx+XCHAG4yPPWJUem5p7kIwL+a0kHXsYnRZIYY
77BfrfQ9C9PmQdRp/Mc6K9PMBGHcYq6RodR0Brm9L67RwdGY54cx9sotYMXLH4sI
qskbtz7gvdN+vI8QWOHFx53ap4tRjO0uYxGBHl1zEVmN7SoPFchRjig2KwQspTAF
7cJWac1w7FjyJAmcfz1LsavMjfXqaYSWRfWRnCjxbP+S8AHBx9JNvgegmRYS2UQI
BGCpYyr8/beAcdSaY1TXTXpLC8J5S+POtBzToslVLEd7NSeqpCiOKPoeNDsRsk8y
O3yHr3rtrfpShZH5IDQCT1U7VOSfjR/1BEQxTXN5e8dtN5wHYbBGtoiO3yZKGPiX
HPPTUJmI093JAdoL9DuGF6ErLJ/uocBS5IE0C+KIVjERMA6sqxQUfsiJg/cqzClc
ILds7Pw45K4ceOx62cD4YtwD+koLyQeRdJnhX9GzPO5akjzvGzsKizArY1+TPXsD
U317Fufq7BQWpFcU9o4kaZ81CguRQwIYezHU1kKmAfR7xvMNKF6A2QTY2a+xh8JI
1okp2NOJUyqx6hO0KBQ/JnQNwOUpa25rvZGzVvMj9+ZbGodr/uW6+ymXzsYSzFxm
XbF6HFvFQYfUCZNVt0SEgPQBilAt1iWjKH2BV+n6g8jEfefkAC1XoKtPxo+jVGsW
s2DXWsc6M5EVQNmN1kJQ/7nNmfI3pKkdn/NB/VCaigAH1UHjE2zt73E1zji8KBfL
4iladf6rUWIqubd8gbiqIqHieGjKY3L33Y6Dol6/XtFbw9ibnh1qOFlKrdSmldlD
oJjh3+3lbedXua3k9k5l9joieOz+qQAzX341zX1ZYUvSoFJY4iX1l9r25La5304m
c8SxbnCrABxlyHFZmHEaFvZ66FRmmdIpI2/eExFG2fiB9FLVGJKvfI6f7vj8EIma
pHVkrauVvPHEuGgEpz0/PsIB+e2f4tFbp3EpE+fI/77qVKh1ZVrL2AclkDTlic+q
hP79ismdIa/kf0b/o9azE8N6LzFyzkMedm9gdNLNrmZRDqS+CRaul50QDvdLV0Bn
6by+V7N4w4y8djslSRtrGg/cEh99Aqj1nnCNYBP7/wRh4ibBrx5fv5xZzCuNsTaz
oJ+3s66iRUXYhz3ayh5w9wLMuc03UXSrKpyGsjW+et1yEomJbfgSq4rDoJoPnZ28
Fe/RoQzcpmENMFX9j/Fs7wWARaZCd7/+GivZbHVqdMuzdsFc985eunOfqVCuOVIm
QkU2JrXDs4Ibae2pcc6mZ83X64pPJ0VvY+CUu4ybcBgm/tmQSdZnGOP2bEgd7R2/
xtsfbHgaRvZ2WCS0TwGvB4KiS/ox8/jsAkvEJbhQVnNLyFXs0yOyBk/pMkwuvKzA
MuFuceOxicS8ZNENNh0IoNLQ6V2I9Sq7uvyDiY9ilwK2BufycZraC3t0seU0ugPa
qQtXbqQzxoR4/AIFhuU5cT1S0kxayZmq5S1+U+uT4YbkR9pcN4T7oKUkQ6h/uNxs
lgD2v/JAhPK6Zf67XYyaPpFxEhviRcFCZTv+19LK3KM1n94Mzj278O0cG04i9SmB
1KaOH1O9bnCHG9pOaYC1wCp1JqZug53Zo55EbngHQQezY5f4swhc3NDqaPIC2yqy
Psoa2Ds2Dk9VF8p6Nipy+PAvNxDqx8L3fZDZxU5HIo/PHWQX9V0WubP73LY9c34W
X/E4ahxqm86cbJcG0rhovj8qj0MKYknNvVHlbH+sCaDXs1UB67bMtOJAt3ios0K4
y6TRqDClDq2ZQ2juqfx9Z2MrKmgAMyhxXmc+N+ek534nQTfs1jVm8SOXK6lIRDkA
ALnprkE/Ng6SK0cuq+oCaYq4MFc5lMZ9flBdeYlgJIKXkyFiUKNGHx8fWw+Jwvo8
Mpf6u5tysUwMmaf00ju231bu1INrKi5FBdaPDJ6ejK+kmC2BEk5H1iDMiJyssLmC
9JTK3vrQm9P0WxixmkjhNgXQnq7x4s3oeQUHV9g7giKQCfG5WRCoS03o2/pvPtKn
eMM4c3GU2IJIKgmhlCa1oXc4KHzpL4rjPI2ukE3y1AcDMgVjzY4h4imLKE4bf4vQ
zSsY0hwXsBGy230elrEkCDQ7qeBCgcUVICWJ67ck8rys0G1D5ezrDn5vwEtDG8ag
yulzcCpevzLoHbrjgfNVNzOCKh+kDwhL/a1aEXHh7Ea0R0PW9ImYNlnn4/2QViaK
ozig2DPh9e9IgDhJwOx/HsHoL/IDI0fnn/2fx2gUNRXr3cPoAkoQp8yGOKYrHa4O
qe7bxLy2uWLrnP3DL5vHQz+R5ANJp9ngDgrpR9zMdkBzMy1ffv+vevs8ofYtfoK9
jWsCrWqO5AgTm1Bz/z8XnLMU1MxJXKS/wunEhOJ/kbElkhD1oCYqfxj4PGlE2OQY
bswSsFRtAQS8qY82eoeK6ZObc+NKbGFXDGS3HDlM1OOxaIqtmCGCO310C8lDUGjf
XO67CSbCvFl7JLVHZUamMgbQP7//xOz1BQptYsfm+fHfPYVM8SCutBbRx8REf6+s
dvO34WkHeY0o4dCF2/E0IFR4vIgOwBKZyVhhuP1lmi5BxB01KgfdkOVeaiyTZzeC
B/9Oe76h7D4DPHnKbfMHuoRVHUoUTpwhW3kPP19BJEIETmFNdveNwqjFi3qmTrJf
0Adrdn6LQIUmCvdWyrc5Kip7xHXX3GR6/3GL8zzGcsLshvBBLsswMKaE6+5Xyfvb
YGn7+MVEKNtS37kfKC4vl+S6m6zKKlnRaftHXTv5v7iAzbbFK8y89xmNB8DuusBE
UQE4ODoneRaIdnhIA2Lk78tXLobF4HLKT8d2Bxl9S11dEGrhg7ZRiC37GoiqoTg/
xsccFjCV1s56DVH48g4c6C8W6k8J/ovG2TJF6lGO4YEPisIuCq91r9CmLB+S0efP
i9llujXYrbKAKPgsV1066Am/p7FlSpHJOXDX1SdOjgukn48T8s4hb83TxO7MK23+
eu5IbbB0g3Nj3SjXlGMN7S6uVqK8J//QPkUD62UV2x0n1mY36vUIHd8wXiofA11e
SFw4OhR9ZN1B40Q6A9OEiX3s1NaXmSceX9uFnHUjsgmzP2zRTscAfrTG6JYRhDgj
AMuWSJLyHfq8hLGyUjTefyzpHKy638uVHY4m5WPIH/uxYra1zGEgp7IvEFj32Q7b
5yqvc4WLTAEa/3hg/8z4hD58RmzEwwNjzCwyEakGu4v1fTnOGVq9a0wF8VFoBxjS
ymheLY8Ddek7J5n3EuSBei+MbhI3KLaw4M2b/Q2c4qcRWIIwq6idqhgv5v6CQkzR
o61yBX8Yvv0iNSAk94+8hStLlNAQJjFi579ay6cH2J2zp27UebLPAyPl4Kuj5BI7
UZMIm+eDhpbdD2IyvxGS2WwrayFOfPg1MoqLeQSgL/6qgkV/BTOQjFGOeO6M5MC7
iuqbCacyxxRKKapIc6tpV2E4cXNq9juaVWJL3AMtB7GOgNRen/TlhDasC487wejH
tpAqJ+vDJhyjdvH6bUoVvmqZxc48uk9drIJKlm2eyA1K6AgQ+PMo0fdX4BUQ5MNe
lIGO0Gu8HlAwHRzOG7W0L7mzqzyBGEHmlo0R0qesRb4OsQu8lWf6J0WxNSf2qOLk
+FcMfGjgX3Wy0JcJ/8AOUO/tl2BaYima8YrYhq1TsblDLm4BA7jnU2TYVvu3fL+j
qyeCCOwUvDU9MId2bYd004RydApmNYNiCi1D76PiOkSzYv5NsFxrVBb+4ltdZCZN
bkurnpfaX7v8u5i/VpJolr2Rb+kSxFyw+KBBRPqq74tXH0t2FK531zEH2aq716lX
ddzs2JCuVtcZuYk5aet5nILLzW8yQC8rlEgqin1bGZ16DU7C8Mf6UZhckben6u2t
Q5ZtAT+YR5BC0/V56iIdNDJvSfaHB4nhMaWYwj70Pwp9BL7/gmKhuHXqeFI05qmJ
1q4f1sZaeD7V2Sy7HdT0CRjHs5rl7yi5gFRsf0uKnyoeP9O5DOgtMRxo6GI2l8Zh
q7GygWf/B+edmtdsS7mveeSc8jD6WJjBigiP7RXThsFFmyOqSBx6Nfmu6aFaACPj
vRw+MQGzdHPsmzMfw5pzMO5kf22qWnAeO2XHxrw6T8+a5FzqSKv3RRpFYBxVuf0b
QlFTvEgsDilbUmmUrq6LEvvOG+HS0mhFzP/9jtETF3kYRHM5DFp3IioSEbsHZPwc
7vTtfeuY4gyiS4R3JOQeZm/qYhLYP+ieXt4YclcjgY1EqmqBDOgGFgYKzm2VwiAL
NrXIlSl3w5V/bFPIb2LNmuPqrDCkki1gUH6pAjhrHFdPrW4+hVDsBAj02KMEDWxs
1y8RfSjwl0I9dRsfeQu/43XfQeJHUdsjMjRgUAeno/yvbiBWsvyvOKt622O6rx/F
LSG79m95txZQ5NArAS+gboMajQx9ugRqxuutby8HjCoOEOT9R1D5IKIxYKryFZ40
vB2Oa7ROz0euohmvygcfGGYsKSWtTpsPCOw5uQ+L8AIWxUksdDpGm87Uiy/aJlBM
+fBqeHVaWve8rIj4mtm22hBDbiLq+gN7sdt1R8mYmIc4ZrcL44ZiKIRXnAf6oym1
6uGs+4Gx94hbuQNWe3AiAUHTlxpfDF2r5JCmAu9eL39+fRSMkHcuMxwDlCCe9ykU
9rdDaSza5ao3itEu0EVYqYVANRPWJPvQV747vDdg7iZX4Nbp6dBPlevFp1vs6261
K3lXarxq64rldscRiOlaWiMIm+1q/+BODZ1KGMwQnB5ZN978j4GVf3XTK0VW+k6U
FAzbYnrhZ21Qzz3ibYrBoTD53yImd77XRU6nX0WD9xQMUUrm7JTtE3tcYdEXi1ju
Sh++1Q0DrlTbWAzweVb618JSc43peyIakvN1A8nhCBWYOghX69XvqH8u4LXrBBrT
MlmeFIWfLxcbs/9tv02keo6Bu2K8J6ZKa0nr6EoYjlieM9iSBW0MF2rnwZyHQje8
OkgyY3o94VEXfIGucbylxVr2qh9zDXdCs0JB/l2a26+r4Eq5vktmE6kjfgVkac1X
whtv7ZQV/N8zrsfgggoxoilDI17dXxHfu/MPLEKMtnZVB91tbXwTho2BBPqbq28t
xsCG4KiPoCL81n+NJoHe6niTXYr5NwNLUTJL4a/BuuL2mcDb2zg/h8RE9IEC0Z/+
yqjp7a9U+T/1eJ1jIrAq0ZTlmLeS4YURYUYYPhzi7htr+GHKnbNTr3UD4P0lQWZh
GL9C2bDfSJvExU9RP34/54ljBzkI4trzTyAdS3hus+hEy1wE4HoVUItpCu3iDzZM
a4txSfksB1f0BTewY18Yp4ZzCyp9k4ym7e7m7lTwGJ4HWbqQG2YXrNYL5hF2k2DK
NmRYgonUMrk8vmlFFvW7NN/22qtYRQRMnKuPO+KXWd9xoCyv0ddED+blz2c1MHHh
8kuqQ0aZsyRRPBXrEUbb88TSZSbDIjlhmvfW6UX7qQZcsoavAb7oVZ96Nl7xzIWr
CgsHYvx+jbylQcw6Kr3cxssFeuw7f6rOfU8nmlGdM4gR6P5CM2IBOW7kDqi9xrm9
o2/MW6CDdPlC8OdjqmVzvj6fsFb8PIk8UtoiJu9Ia/ErngAL56/jqq7ElFe9zrmJ
+s0H52U7VRE8zBP51W1xH6CC4ps4JzJ0Tb5TKS5yy7XvxDh1WGWwJ7nnwUCyneY/
c0E9auUWASRBbRg5xEyEplA0WhscNq3zRF2eChQuFzpDwj7vVuURodvbv40IJnL0
lcXep2mzvZ0AjgKXkdDYyiC+ytMtgeyZ/6MpXZAm3lg99ZIdw6JVuchILqiZPHaz
jbLcDU+l1eEnlUGr4vusTYv+2yPrgQ+f7QWgn0nCRsTKxDunYk/GBH3526gbq5vp
tmhkMlUEI01m2x9FPJKj53PHwY1y+eASTb5I+5fPqCnFZdV+J6Nj31RMi824sz9t
zk1qHQ9Mvtl+g7ngz9rILTsU3gGYcR13LI4CbqUcnHPLXvN4dZxHP+KMbAqRwg77
6il0ewU+UoPqraXQYCFe6wooi7/Df4NNdvDxAgoOy5KGIkKAWCCC11tLxIhUFdtz
0hkBAnMcVvRx5r2NpY4Hpc21TsLvG9hl19d8p6NxkPeBCLH/NUe3ja5lOS7lMCye
Kvq/79dOg7hwhjWbuNVQxizD4BCri/6AksEBSxe6qtEGR+FHqtjbCsq2GNFNFLnF
sFpyfRn888rIiCd4dgWVjYx85gDKI9vf255MLXmJjUUGMT/ptXe86PacvYs/69qq
OfietIUYO/vULJhhxoc7e9spQBdpdv9aR5lBK5JWx61khRlThOJn8tZmc116ADZh
tRH0NX9bFSB9ytcC1esklcfhwcrzqd76YaKrwE/PoxcvCnUkpw2PhwEvdHIMW4rK
7FVmUWWCDAzlyPxcGQbTtV+mYrEegNPzqXILKNBTkYN4F619g5LWVBXygCbgq7qv
XbSHdgEqpfwrPjDyK68emHBcCPaDEmRML1AjBMaFJJk/0Q/iNR3jRzxCfLsCfEb5
2KDghtmcMXQiHabS2mnWzZ4bWctoZFePPuzs0pTDggIOtpimbzrr2i6PYOUjWg3m
DVB8bSsjrDthrRcna8YhGyYn0VxVoxDgMeKNTGO1UgxpulsHIisVN8b8WG190M46
zRRVMB0vY9vCP3HtC1GxXOHUXgL/lfOx8d8bXECPuwg9RO9k+PbNVRcbUVoh2CIr
knFqytWv5d91DxvK/lc3Ug70aKozJG2Tj4R1L1FmV29hy0h6iq/rZsByOGKbG7+3
aXyYA47pVkGrnkROrVtgL+ctThwegF6tflVHUFmJuatct5DYDNvgWTmMF+F5wDmI
b9EwysyoPW4OPDL/o44R7ygsvb03b94RYFif9rtUlvqT2YYYoexJy+TCGN5ymiQo
fGfkL58JDUcfpfWEMzoCHy3okdTDqSwG32LfkWRsf1ojqOrDzWr3pgP4hNW2edjQ
dO+M4rabXCOXbWK6CJZ1335rf2BZNlABmqbT/xrWyQ8CUB2N1Sw6Bw9qa7KlC6LE
fqLGLDhbCHutBs4xHvYliMr4EYCpJgx3uB9/DJBNFdEvRRhA0GrRqlBattzwX5xQ
EWB5H4BN8vj9yn90I0kgXS9pkZ6D3pSoviPqaJ56mVqbQuyL+y/IY+EoY4kZjUpW
EwFygTD86kpeEpAssyh+15wSu6AC9NUQQsY9DrrwC+80K+MwJhyfllKBxa6NKwaz
SbxfgjASoSoedr4nmhwW1JBRskPGluQv/6EZ2e8xi2dfDVG3QA9K+5LZjPR4/vnk
RPKH+cGiXGnourWm+sRQGoHv4AYuL02Q0HLmJ3K+ILW694PecYFjpHIdULHOxQKR
I/QoYZ0CHHOjndfxNjPOhARoCTSsO1e9tbd/Si09L/EPK7nHf25h2WxA9yjjw3PM
u6e1LmhQSOlwqmgtQcyqJnyvpT+2o/osgxN74pWuSH+ArhCQ7QQKe7sUS+9btBgd
4xTDSq8rnCZpRWveRNbBMVRetG2h3Ayr4QQnMuyDDaacMI2YChD7ZwRy4QH2+poy
ROMQI4eUJaPm/wXFILEQT3axu/ySHGdJLxUF82yFOO8asdxJhW34kwY+eIOE+94B
PYmMtKZQhhuprcNZm6pmWooAaQDaI7GbigRvDvD6MCpYFz3s4XOdgyrctSmhHpIh
sh8DGgNYMm5glQsHwk7b3dfrwH+q9/aOuMp1Azcygi3S1XyCqsr10IvhjsGJqk1d
5tuVYDnMSqcVJK6sw2bb+0PBn/L6jdEDoCy1M49dlIzP5/oPdUijpzeEptzJNZZN
dmjjGCsB5aO2EpQdBm4ToSZZskeknmOTqNDjdYfMaJjlfyAAiSmUICrDhJYuWJJj
LArSUVtUOmeYaUcjc75TO5gb6DBHEf//JM4SecFBQ4F1CwWSQE43wBjJgGOt8lSh
zFVt5mKBifK1/vK8fHMa0aapW88yz3mNreNVfVLHHDArLANwsjDPg8G68liHyg2y
G329C8VtsPPokjHmHyxvfoBL8l8cLiBb3fLvJmTzR1PIEqFHy8kvcamVjg/41MPG
ByfziRt9bOKIHUCu6Qw9ImAZ5+P7r/xrTZtcDoU9RT2aooonUYm7vxLirqBlKi1r
9/5QrMRyVhYuV1yaTfxxhza7k/jYbSsaqTjIcInGRNVDJj1T1ODgFfzKkU7kxdbZ
pjpJrUfLv1p1gF6RCd0vVzafNa5trjie90cwNDZiqpzrjOKdbfR8y4C/pMoyrXPm
Qfmmn9K13C8d+jRgDEXfhMowYx5CazHifDOuFT6dcO91+9oCrd07oKMQn59wH3rs
wjZolECMQemaE1sQYyh77IDTChUM0wP27YF8dCNsYmRfVeb47a2s0SS1vqKLiRUp
UKq79sV/+/u1LJHv9Aqq7cMHqPWa9XzTq7Oztsup9SnUPAag+IX8+mzdtcMf7EDa
+2ovBPwtpDRWPZJEEYPB3oWUxRrmZkGEkeNLsrRc6+f6RDfMFmYem3NBE6FJHWhi
iHJEhwxAX1no++qaNlzuCYDOfQ630pFEwa3gv2/HmquROTRp1vSHL0l5xyIpRRVQ
n/DnNNCaRia2TGyIT/mwZXFYETjgDLRgHdYIQu2yVU3H1euXhxDcOCj+N/r6/YpU
RMV9XAfKQeqc+TKGAnpjuwFKvu7ApqAyuYsORxsEoLVXjeg15rIwXbAXHTpSJipj
zf8wRsHj5hbjAEA98kVt2XShW6fq611uj9OFlR+jWfs3f27xIbJBrOu1lIRYGrvy
pf+SfhsUvPysZkH1+Mg+37gO2dSU0VMR/JZtZfhX1RMIl4qeNmWnvNAVRw3SaNcl
gOYCmPKqQn5GMiON8d/BHhdB4J1PUEmVcqfJMoq13xIuabYj4kHNceM1QFZpDMGh
LdTPuWU6jAOdkR4Y0TWqH1wKRLnBnihzDenafBbhxMTHK4tH+5mwFdw/euvCp7iT
z8uV87yEygqP2OfvD4KqIBZyMPw02hju7VPUFgTxicjiEZAMwGZGoqb4rIxj8kD5
g18jci8PQ5vIlWZMeIQPSEgoUAhAQuq1/elJQjda/EKeWirOkKMxtWT183lL+d2V
vHrp0sbn55z09ji4TVxM2odp7zRF8GzB/tgweKaNrewEyXDoC80zWdV7y/x13kXW
B0AXdsaGQWFnqlfWvq8ZG3UtMQju9E9XwQWBnvafMOf542xFWND0J14Zyt/dImLk
hAfkUIelOREATJtqWecTFR2YdauNb6hdeGVaoP+7dgtmUTF4DXbE0gj8kgkxy//r
NQsYX9figpeuOJul4EAE+FBZxwtieN16W18JCxCxUKull191t4QRmSQS2YgSMeI2
RxY4vL49CoW0gxc30+5+paK3Gr0F8ELE+eCOqYmYKV5I8yoOcJHxEIH6V5Ym9R4A
FYqIiTXRDN5uI9DPdoC9FL4lxyHDHr0tPZng5IWOah81jJbdOTt02zbHLiDZU23v
C0hu2Efe/7C9++xYCMVhNqu/+BSLfo0xwpPb2w1LmAix3p8TV6XFr5kncU2cEOO9
/fdRfvK0zVSq5Ry4FRy7kb2daWx/ndKzSDp70ST3HktLIe2Q31/ChE2tTb8O2OAL
ladoCe7Jb67Knb/YKyXRm2tVGhDqUegdBTuM6W3QlaPsA3arx+lBJYjaHKvfeb0K
c8j11EcFuYuzHkII1U+ttJu2krrA4QReaWmzxun/eOy3eH4bqkhwEgpeoL8QV688
LuP2y/Tu0Yjeef+pcvdgmOYkTU5FCFREbtMoZFcF6y4VDGASmzBlly2T4ZUufXcv
CvdRwiHR6nt0RcCqckGRvtPmx1t8nknNAQpINX1wpEK6R8VPmiG+BZlG20G4Gp+8
UHx0qjrPbIQdXTUQFlUHfoBx4niDr6iT/pWoD0Exv6iuEtOmoTAn8eRV7Fke5TzP
fbTtPbf82TVG/BVQZJQL92dHW9nuFZNfrdm+nNJW4Ys4JE86owr96zxUm9WZjD0P
zAZMWtRB90+d2aY8LQlce+71vWw95y2JtCfMzVUIyUzJ+kHbUJsNAWXn9MdVksfc
CNesaSjGn9/FdR513LnxnYKXTeoR8892fBsOwkB+p76yqHAVGswgw5/KEMvJKyEB
wLK39LVbMUAC7HLEnYl8g8mTN/F0rxK1p/6/x+FC15ovXMe/79TEWdP7eV3bCdGv
bO0RvFh/UU3C8Dj2f4UxFIKY98sX/ai5eHaNkYiV0VVIDBKkZ6cFMsScypib70bs
A6hUZVPKksWg7iuAhsyleM9EFR2Vv59L75sa4trmyqJ49zAxZbn1743yiY89WK1w
wp2+KPsmODyT/riPTpOyC9q5yq/S+MYCVMsdD/PnbczCuhhgHMf/a76WhB5GB17Y
4zuVK1c6wZkcAiO9n8AaJdxqIfiEBk5rtWIH5dzpjJxTlahe3OqQR66VGp1knCPx
mJu2kN2kMctnwC1lvqhU/wz0U5lkf+uSK6T5Ws0kt05/49RbSvIHNc7zaANSVjRK
d2YmieOnOnqCMR7j/4/kuARnDq4sZdyCEreuRUMxHYDpai+b68YG/ZWPVFG7ToOs
FQAlCuSy42CrfXAVN3FKiabD1fq1m8kq8a77QG2luyEL5pV0BA6ZZL7MgtkePB4p
a+Vj8L2GSNajx4yUei1wGFoyZknU++OXPkbZBUXBq4BrvBJ7x64rDOJNPHSWu4p9
W8j4AXa7rKRxXsx0kZEVr8GH4KdZ+QsICpC8eitWxt7m+B8N93LK2AkrjKGUjedF
Bp0fScshIctL3iUYYb6TVFswgD1oKzMUUeNL32BAKhyz6KANuwqftNEu6n1qO9xV
B2nAC5R4ubsMYMMPDH7VhlosSENhTVRJ9xdNH9+LKSM3hiIUAIDydBbKbagX68F/
BRkoutC5Td9J6rzqXcWq67mBYs0U0OCuej+Z6NC/KWHiLN3UlBB3u9DpIlyaMtGC
ouTZPLyxKi6dDXkxgqjh/6DrAqEPeJgbr+LdUSbAsD+niYRq5zUr6yWNR71vMAJE
uk0dsN9Je0DB7NPzdlPBSwAPE0K8Z1zrZeaG5mYhhq8MVryP2iPflBOP1OCivaC8
X9Jb0DhB+CdHENdvDLaFJmxdnCreGHQvKgaGtyP1JeFzLG56V/J/8al05nqn9GWz
bbBZABZSCA/ezWvyyYlWw2fUaK/rudg1gggIbaR3mz4GENS8Nq7DDSosLK12YnDp
v4CwLJUQws0PT0ga74oyVb0EjT2CU0v6GhvWV611k+FLFS7mQw9T7u2Ey+Yc5q1f
nmNtWHO19MUSKQDQzlaCKoHawGAWeP67+agTOQzhLGxuo0cVMu0hsj4JI8rp3hns
YlP3Ajf6xdP5tERDb7OfqDjtA5fBNaol1E+7DdH2FL72oe8mWHzvpOZcOZPwQAXI
3pWcqI0hj+05RcQwWNexGR35ROb2RoVENFkHK3ehIn6KgPG1sBhdxdUL5i6JwLY/
/I+ZsXE4NSItbXOQzT5FikU6gaMvjVWO1GC0L6vZOOgE4NUyzL0YFUma2Z2OkETd
WR4hT0CH/B8cCg7fFdix6dA7gmZImfU0028LBRRTFWfiNjARd6UqdaYNxqOxhc+0
WpyzACle/NzsPRz3otsbwugCGcf4bKh66ov+00thC3tCG5TglO3R6jUsQFSmbMEe
gC9orTWWrWd3UiDp0Q5Nf67RAzFoPRd5dL4avHNp4qZboIb5nFFfNAh81WvtorGA
8wDhyeDqes+aurmuefNNIp0wCGr7iNlg38uW8E3v389RDmlrD7SoWdQvZsSglwN3
zx+/EwI1asJYt21RnYTkuFnjJ0xMozMbt40Id6M5osDoXklfxnJ2IXo0d5nSWc6r
zUQHW+7OSxB1RRoQji7rtO5sqUy3KWsSufxq4jtbvbAy3MpCYlEIiseTA9HZyDiL
J360+wuSPQm/p0vU92uH+TY2nyb5OqSFdaU4MXUrWLqvclLySsaZRmEWCd2YYfL8
QcNDa2TPcHECTEeXYDqD+IJhBHqIK3kOfnr1mZraQL8wY0nL5MqwJVUJRPmFn34P
Mn3VFwMcfZJQjrXr7XTdP4z1sj5RhrtPngUNn8GlYfEZOviJNmNast21iNAxN58J
8xQ6CPt0Z6NusjlB7BysVGFfiq31w3MqbSk3SSrO9oeo05IVMUmLhIaMYNI+B4Bs
hEoSmgf1Rq/oMrtJVcw50t4gP/3FEWbJEdKKzKFg+JFsNnasMztP2SFdakbQNpvC
SnWW+vaBTobihpkTrtiNlXPvE+Jo2ofw0xf71nypFiRpYRclNMIme0YFEnv2fl2o
MaRGXhLpWGa5BbzRkilPBa9p7m/cDkvnTjFEwmVbrZZhRIBIK5VZ73s45kczD6ay
hEtehxIWFyVwM0XJFGPQh9uj5PI7nCRS/L9EYIDwvxvJOfD8Nwbh7mIR8+q9YBD1
mQvcVlvoI+zVobAfroUunsIQZNsltf8bYNlsph66Yda2EeM0Iq7W1iE5oJGEKQso
Wt4VmbUwXAgN580fFPruUx7Kd5BnYdhlGqHrXl0/d/rPyFR/vbaIzPqSA5H9SZyl
2nb7oQBxi0arVOOLgvc6k7cCzkcC3Qo9dEdT2t7689IN6NEbsAP+rsfD8GTNt0sO
tENY+HzvTHWEiF8j+eerQWMwCKjkkRXzF2x5ZFcmjTJviDXOOcTF6hZ4UlRWWy3s
45lwzggRsJD3LOZQqJBUL0zNdCgdpPDJYLLw6NkyQd8V4exlmVmg8ds5wtXUCHY7
/4Fkol+Kf7J6BEJ/buL3ul+JKfdlmNfSbn/2CYkGX//Ih4CIZuc8LXqoKFOWJkaq
rxVKQ5ACDRV4vyvObDUXK3GFsz4Jgw/xXHXKjjRyo+eTOh+yS1GXXHwHgR99UfSk
pju8vbw2YznihnMQ3xkED9NJfiWVxRtImShbrHZIVmC0aRqNhWsCRjp80gZXEiqQ
Lfp4lAHmUBEw5EaMYVZIVXjePBA1mknLa+V0vGEPVPHuAX2kadOIeSVw41tXf21t
bmMiVfzjPidhB/t8tJY6k5ZkpDKYKioeo3JnWswc9+m5Nrr6lLNDOHlVB/5f/60x
TDZFKgA55vZpoH55Y3qzPD6Was0xkvWZIxeSq01fZCOlmBVRXKTdTqvLtENBkA1o
bSYmJD3xIOvIL8AT8JjSC7di+Druw8xn4Pj+yrAzq1tTh7EOxbHrfXcmURQxZjzy
Z0/xUVkkNiT5g/iRyExW3URPZ/iLHVOLMbwynwsHwtSzVkaR/yYzZwZvXRL0qIcH
DaWPckHBCUmAj8aZUBf8dBaU2xi+mR0vD4/Z+kGVyPpF96M6uFwFGXF2NDB4iJMx
wQrcEtv2TJVlSE+omhkeEStjvqftxSTOqjdBscmJWe92FzWNwpgtpjTdCPwUQ/9/
eH9MEpeJuJzNZC0Kc4mtAORv90PSnpGHPXyT82yj3Q8/u0vXTKBnNpYPdAUq+pT5
EwCTkrs7bVZ8ImMzsveNoEa5//IhwJNL6u72aaNy++r2fccF38/bRCWcnuPtFA1U
FaTE39YTDf0W1TsyctMdavLMRvTutE35CwGU+NB6fhW5QvJhxvvQrE/AyCXtLPGm
DlELivF/O8MNriSRp1ZJum8NbNCjOs6mpbWae+mggu2laJxCy/8hLl3YgmeKp7RN
0xVhTRQ0Dzr9GEQJWkeROn0cYyRJBGeALjJN75yUTMY8wkpZ46Ke7uRLfzl+OLnq
qsQAru8Kj4Di1wmPwGIyEq8nolhZ8VilnZPXGQUg3XvbH7oaIoBQeE/IbJp9aW2W
P7jsCXHr3Zr3eFT7IeY0TDk4OlJOUFOH5QSlyzEfaFOOar1d+h8YMHQP8a+/OnF7
F7ED4FW+1dUubFxlcH4wDvQL4K2nPdvlb4fdJmVk70RcaV5UoQMY2HAILAKurcrA
SsKnYPqDTGqiqgBCEXGFUCym4JcFIW886coCHYwFOv6pLaJGmiB4iccziO+85t9B
ExlhQUv2VEbzsc4LKDWHQEvTO0jnUmH87T8MJqpLNRlI6W3nu/+toRrMDpvmVePF
1uOt03TWypdzB8NF1vXp1TreKMLpKE9bhohI63LaVNl4bQoMmfzm2FVM2A47caDL
hp9RlB6Mg2ksAeIEdJMVXeN+NJt3EJSmx8llZIAe5Yv7exJ62/+YVKV50mUX3c2e
pkHtTWNXdX7BDKfrNNoEPQv/3/lT18E/Ato8+hBva7CA6NcmESO/QQ/MloYCDJNl
8MPLpdyWm+T40lxWzsFqSB/asUZbDVlb4EbP2rWcBA8bgBuFcriSuu3DMCTLj0v8
y74f7JNWgsDmxDhBSzxboZn2iCvqD12IBNto/2oRNJl85gWVxMDrCFtay0+A8ISu
O7besUe6nh1zs8gGQJWtBz1wy/j39WzqkXGjasQhVhhjgF5PSI0Yn/NUUuYwid3L
zETG07m0VzdmPNuihTlIjh+mKtvTv66cmbUzN2DA4auvwUknvAwSxpqCf1QqQUZO
a2xWkm6n4Nq3G9OnXHIg/jmOWUrB4dyAALDALiGdds+Ba9mlRTrieG76h+QOOmtA
f/gFOKCkscKKjDOz3EschXDi0DyjjQvTc2sN6malT5VJr/e/SUghcZrO5kNpxohN
jYDEkLynVdgfiqqoEEMrpsFez5hTajjBTA2gtolLdh4PimTd5TXC1C3028bBo3PI
Gto243ot3BzSGoqludTlEyKfIXqEtxqg2a/LSDNeSByC7p2wdzWIvofeV124GedQ
4wa8+61otHbYer+XGxEL+GqEOioUkci4AQ2akpe+LI4FzJP7yrvx4u+ofNFGbArY
pjjCm8I5YEmHIAK1wqXXP4m9ZSvfMInpb6R8AKcw9sOR0wiH4NVxdqRIyE6dmzBF
sx5FAfTnrvuxpa0xDlLlkOyJBVNEXD/UpfiG/yewxB+qOsU6ipRS0wrNiqN3xG+G
c0LGvf7f/5Yjr42SXrM6xXSgX7vPC/RCFFqQg0qP0pQtaU498E8BReQ9TvnjnvyD
gBsI1xI86fshKUwtvkQT6WQfSczfMiqTHs/xYDuvXUpW0Y8N3ALPP7h+j4vo8nl2
VEoQcuhpeOo5PLNpkRaX4/KYEKMRkEzpaa8Es1A6B6tAqDCesNbEBCM/v9bap5X3
dycjohR0of4isQyvN0CBPEaCxXWAsVqR7C4B0x8q1ylHkt6R0z+QmHvBg4pySo0D
tNDJPbrRnx8tMgv938aZdHEEunENlc91c/JWs4KOlwz5UaYecaBLkoGxiIzuoGVA
tVvWxbiVnL385BD0AjBEEtnWlNtO/d+vc+qDDDBQmHBsgOSAtCBUKMZP6jsUDFii
dB/+ygUjsWOcsycTtBRwXv8JITbzntrG58lM8QULoDWSa5flJyIt1+7Mj0Jdb3Kw
PuU45jAAxXtpoVHzRfSwDieq8DTzaytXct09ONlJVGdouAG+nXNaJZxVfKd6NUxH
U1454BOri2fKDtoJt1KtYXaydKx4uxryd3PNUaXlPSW+GDtphkFbDNgLYqEpEJlu
7HfoLEjKt0C9QnI0xfEH253nYgZyY1lT/IDlgIZb0bC6bFujbvdDn2K10pxmzsde
D5Qbe8CGzGhaOW3alUR4nw0SVfYmwf1TGpRGN3yqhT+5I0nfv3jsTWe/HFP7hTBT
F+Ru8Ixy3bvtrfV/A1NlQRi/G8GitkbHZ3qn4ECyJFC5jTEavWzN4YClctcq1ndM
EvzEDNzoveiCHWrfRgziA4H+CmzRQ8Tmf8k2u0yOhLgID2E/tv9i4l79DUxlopMf
hqkyE47CoTZpmI2yZBgzeLxpJ5JYdlwwlhHVqUfDwyoqfNx5+9Ts6e4Aw5kE8hxP
GqW8VCUFDq+JYNKnKKDHdca/PI8zN0+pGYTxJ5V0eeLW2VP+vpUGI0QITD1lFHwh
YJ8vpBp17xwDhnEL5OYzkNw+s1daHWD5HQHSZA6u+/cw9DJ1Ij0kjfrXwdPFplom
qlH5Ql+QwVI3Qjw0bCavuOzWBp0AjJQHePt6vbzmHIDvycs2N2DBEo8H/uQEGmJ2
hkRa1zfLW/S/SqettkeSvDoJTAX0wqYdXUT6QC/RKRIlWDTEAWIvixKhX0Ufa/qD
llZeMo7P0CNziL6vxfx8rMotXaMosd1ZIlYWF7MYQUE5CgLp6apYqO76eCfFe34A
fySJpwek0qpfneKXjlnbACQpXR8YixRGKmYF/U8WY6t2aAG7Upw7F3EDmQmfO6oJ
DhuAdYM9ZpRCOz8SGmydQzhI0ozsMQqUxQF0kOOOD+BijNbTJAZX5WTcsCAzCUGj
wQI1lUcKDDbxmOmYxyP84/Y/i/yxlqgkmDqV89PeNfvZ/6hWUhB9PZmuVIVPjMyf
G1PgJC1S6ocgE28TTrfpaIPkbrSxIah207FSrUe+9VpP19HK8A8jTK3hvlFxjMAC
W9o65JhJ5q2h8IHhYW3XS/WNbZHh0BP5HBRXQdVcS3SKydiMg96T4YzmtHT2D5Jw
oEHx2VhiPBbUngZcfBAlWPD+uSzaXLttrVs5iqjn85Epx5w9KDxJpX35jn9YItrf
/br0J68RC30OR8Bb+eDFGtnZ4pJLg5mchJriHUytwPUtt4n4iWcezjDhhE48mWPI
IF0gVuePxdYi5tQsIWH/ghkU2CPCts+qfIt8AxXPl1HJqanZuQh4N/vMy+kfY/Rw
kkLPHoJtM0oJVXBCD24UJdGC5k07+unc+ntCmmp1sO/egbs5mW8Kymk80whOo/jW
IidnhXLr2vyDLDW3aubyLHaOlEJZlAD1u5F7mAFTYOwl1BvjYY7aSiNorM9GpXd/
94pj1S8o9p31A+a85AW3awPxkhZ78i5D5Eivp2Noz/OiXuiqHedKbNNolj+oCThj
W7HsseLEfTpFghfOXKt/VWrTFneO1oPewcBASkJ5dSRcsRZLAAR/Wg23bij3a5x5
dY3W8UX0h7RIxO2XDnFBGWYKQR+CwdrECOMKbvAcLlh+pEumSkE/+Tl+RUl10KzH
5T5jf+W0fyJwwv5Lo/foyxWqsc39709IYkw1y2M7OO44abIIadmHJPzdaw/uXBJJ
XuG3iZfBc/z+FhK1NHSe26PbljL/EOiyAkncYjbKQQPZuWsmJFPsp39/beqUQDA6
llCeOypDvkPlzTagD7nBkQcy5B8b20NzCXwMOR1Pnbzpvzu+gBijm32W+SBYfIU+
9uwPk+1bcfVSuQ0o8bopGS/nBHxI28U/nKNxXIWS5uyBSgSO2FAa88msCajoeBvs
1/L8FNjFPh7oTNaod6rpDfuTJLjXKQDn1cMNFTjR1++RHwsZaGYTfbfQ7rfsYIiq
N0wVuFt1jJ6hpEgf3P1rYV+vmw68evQk4YjhUTYlZuHEi6wYJKzOptWNkCu+xbDX
v3ovqZ+VdA/GOcB3fnPkHVlJmJVQ6mRfvINOCA4G3eqAvTdxGZGuVWiKbQNwBWoj
3duFxJ3aMjOuxgB8Gr4d1iDn5h3ANOQOSg+LmiRsVtCP1+TEb3jr156LWrbsUSMO
fb1gdGBof+YNshZV7JjijEvpE5RZwEngbwdc/lpc8uLT+TRl9xx6L9lPCDyO1u3c
0Y08O5fNgoOxJz+QwAAgubTGD25+vR92FKHbS/FHIu2BS6CgpkYsARl3JQPOK0t3
p504OCvYz8mrdbw53v0ko9J1hvn7233WlPacahGW/iAUwbxVuLJiLRMONm9X58tL
/AewJNfyGWocxvPMjfpfJNpbQHDSVjGLoaHD2K26WM3sVfDPj7gO4TWCYztkCOAq
KgiejMaaKP9cG6be8bJqaiU51xppV4RsGxRpOxqwFlMRjefnTyJf9DzhivpPx3V8
Wqztz8JpFJgFGYWwz7J0YGin8NlktT4dONfVshH5+U5TwvCyqbByJvESYw8smizj
iMKaLswgf6tNtdCV0YHqKUiad04cyo7Z81LSlKe1dQNdI6k2nw96PIFAimf0UGPk
eNXDbHCXpcNc8E2arzJQBVQpSPMRWwTlJcxuuPOZ5hSX7Zsswkf0oyvmkj4LsumI
0Rto6EQlJ9bw770SmMGADgv23mVoEHisKqv/lkwBPNe6HGGMW+GuFokzePM4wuzR
kJAg6uikGfjHaFXSi4NXEitWK5dUWssUflZdcyddmSY7imbLa7k0Fv8cGAXqFmxQ
c7NqCCNLM3TFufBNoHeHrewj9glUec0frdfD7L7dzr6WZ7jqxw8D3pqznoU5O4KP
+1ZuiPlKW2sCaFI8jdWRQlUcvBZWqu0h6NPmRqpc8znB3M6YM2GmQ8S2yiJMAuej
C1zwHmYW+OybhCUb9gZ7FH79KZPfXXMh2QYkM/iE3r3e2KdsOHjOtW0unBvzkniV
h7Jf9G/trb8UWknXfTSw3y1W8gZu65Lu8gOC3ug6vZ1VWX07qjq1oi93iTaGYFj4
sOWuF/xApMJfMwlDU7hx1cszeG7Va3IE7YvRBDRfcKr0vsgArEUfsCfU2z5NcP6O
vMbQDhwDAa1ewmqMPBItO/SCEZ3LYzy8o2soD3CYOFH8y82JEdjcvFjE63YfUgZ0
BK1zFy78/Hkt8L5y95/TYmaqjVM9TKb2LYYaGv1g3NrD3gJoXBEnrC6xHcnrMdmj
ixBbNUDsFienKPHg+4qvaaSsmXwO5bfE4IQWJAydRMiQtiS9z5EoPwMhBBlALzl1
TRRKxfgiobmri6D1Ypdiu0Y5hMYVyNwD+0dg77IVKYjvAqdJ0HZmC8kv6zxUD8Oc
lhmJg5VcWetavv9wmgUkKh0NOupOz4Nfk+LARZh/rE6+0jDS88Xgz2TVdJQPEfmo
S0/Fz5zCDMQ6jfYK3fzHztrJeEsF2QIrePzXMjO8Ix+TmHy6VA2nah7oRukQ0arU
5Hon9kzzgBeckj7WgL+4GWtO/2fzKc2RezrtT1f9R0kIUPy3qr6KS5HKA6lwQJJO
df5joEYwPD7Ss6KF+b9T8ALYJtEzshE8KoPoFv47g7utRDkgA4KYFBTlFIBzQj3G
3GdJv+IlduEJ1pT/cHlnbmhOkgjys2krgNCEi+NvlSrUwZKxWT/jgq4MICpwcChH
kaUNFHSiZz4QTtSpMcasBnz2gPtKd7p0aLiodEgrXl1+6+1uX7FXBgsaHqlRwzHh
w0o53dZABCKTp6/b3FIYXGz6dtVKi9MBIYmTtRdyRIIclcJ+zYYKHX5brjNoy+C6
EJVgEfGcyTUaFcVCxsbdEnf32bBTmrvFv7SLd+yagwo/islSr92pLwJWsHworm/A
TtweDdvi3I5suJX6NppuwsgLNb96VrnH4R932BVOOh10XCwm1pKcyLvIu8FXQPtj
RbnisxLNyBAFBjy5lLzXUXMh5UKVIso9IOgpkJdjoswiFaX9X+3LO6QK6SJuhlPG
rTSAoeKpjdGodRHV+YROjvJuVL+if9AqUcFH6MidwyinzswiKrqC6p3AJiwqkWN+
W+lio9ePhvHdREsIwPhNnE08pui1xEkmhxSZWkPHAe5FzwMD7SGm26k7RlfNlG5F
1R7s5Sop4PRyEs6lkhj1uTtk5Y0RpX+vqJKcsuW9U4vyzLeJRKBAjbU8iPmsuqRT
Qc5uaw+Xjw0bJIlqWMyN0e5temjqpBjMa/WMv3p3a+zAZS0KFYbuThyZ+5hPweGf
4upm45UYqsPCoIp2ONNY1+e9aXBh786cO8JaHcWVD71RGTeDfh8SI2lB/iG4RJgR
RqU+DTXSwYlE016jCFG8Jj4cngjvATZWYRlVW7ngvsdEYt3vCgZQPl7Vh+MVvGEV
aE2BuO0hUPcvoxHHD3esvNN7VxrjXtiJ1b4hklIui/XQUwg4EBZC/YVyHv2i6kfP
z+0ix1Y6VhjhpbCJSZIF5RH1K02PdzgZ2eyoHCZRApOEZrMTrXsX4v54xJflczne
2rugLbOjtVLN3HuCFFwkCeYJrOXNZA1V7YLZTKfI/85vQUbIn62dW/GRj8Z7ikZS
8bc4tUnKU+Hi7J4zz5j1r9d7FBye/jXTQc6x2hel50MW4uwi87EayIbXJBuzBJql
7xzzn999fZyqz7q98kn77OS8yO6hcPxEM7KmceplhGhf0xWJ9uuqlmJDwtWvZBY4
o3citVNwoUHVv35zlvjT3JH+bVPIVXaWj+UKR1XXeZE4FRDLLBvezz/z0MpOLiE8
j/bkVoTTD80lk1Lj2htyYppgYzDJ6bYL4nN/y97Kci2/nwUCOUywdLnIFSq9P35K
7jmERA+g1ynR10raKGT2EykXW8RQBN1/emPyWGLv91vXgFx/9NZwfyhlKnyNoyui
M8vZy6ypSQJdS+kVe+bz+f1uH5Vd4daNlj9FmRcR07dd63h78qzdddY4MB6j1dDu
Ic67QfqW7I5Mqg9gSVp7hfk1LurPMC5z8YUxMzWw3A+9F193YnWvJRTRY6TxOCbx
k3PS1TjiGjSAtGma9eYyC0b+6y3Rd2Q1FGHuFRwX5ecdP7WkRD26pT7VVOsVAMge
YnIL+ggtWWoTGZ6L2E5zekoOMqFXDFZTFfpLidxFpUxEIIOOWSir2eRIeRwHcYMd
IQryEh3eQNYb7LLFLg0hoHN3gvbKS9HOUJMXd0JIezVVLnjvlrapDPOC40R2XNLX
oQQ5nVxWzvy6S6rlTwHKuo2lxQ7Onwlrd4nqSaD8KSdmZAg7QMOlBgDnfTagwIfO
bVCiBmMYSpxd7OVkcxY78YXVjevO3PaxMI1xuBUXUEeMZkiIJIYrY66Hx9IM4pPC
bxre+CMl80xjzhVAqDOX0WUnwq9RX8jtEtSZG6F01UlnKv8GHoinx7V6LA8Kcp1s
9OyYEOZTSTrhImf7P6Nx0WYwDIgBX2iyTHsbcMVAu1gXbA18NjzjbbZxmOsU8qzV
4puSMtq5JWZGSRdsSRXaKSBGpsCziXqN4RcvE8/XUXbDumJHADJncFUopPWotjgd
tVUpZ86xEJ5gFJroMlYaeGxL0MzpwVeHr5JC+/2WBIKvuQbdYlSP8OC2IiUUOcxJ
yPMrwMhBZ+E6mwwigGeJE1FOpWuXc0VGuLURvCPvolRURojR6C9LVWdUAI5EC0Jv
hDMYOty4NYjsH4HYKD2v/EKdAHJ6u/JNDlM9gjKxS/+8vcjupWBxTA/IoiXOMBVd
IsC68QIurOBlqr7Bl8jjbuJKmaawqjUE0mtm0RpAsI+6GhUGTMbM0Z7YxVGQHCm/
DzK5Uk0SKcWTyO2JkMv+uhKKwdA0xTPolXkXRqCVr+5ZzGXBBsFQM29W2s2bEqoT
rn/7QJA2eLA26Zr94kmMyzHG7JUOwzT8RT866V85XqC/03KD5swJpkfjqgkAba4f
7fOkPKyq3ycMYUluaRSJJpYhReONJ8EgqNRzFyOf9MKbXAqvkxmNyP/pHo9FQquF
iVxREuUj71EYyX1RJr7lg1XOgyZ/bvFXoTQSQieAPCx79eVMTTrrkO3qAPIR7Dus
j/BLT2/ZHmomeszksWsew0sdS9a0J/KL6tcUynK6j4Stiv90Dc2Aur9KsbDtGH46
KEI3jgxx7rYxdbqlx8htOTyWEJkTb+Gjdo+Nt+0q+5amqyGtmXUT/D5Svxuesa7q
S/1L6weIR756Pa1obDjLORQNyQrv4fLhRKAIHDAIDz5i3pa/0EmZ6cV5c/H4hxaO
qKM1coiaiBuf4JnoaX7ch6+o7sKJq7dOKl4t0l8UMA7UmuJZ6VXvrLkYxPXtQcmA
LwAP2bqgOcAkEgl/gMUNKsdzBny44ky7hcU7Ty/21LeRn9crYQ1gH113G7bmhbCx
hZZ/fh/KRfAvtz6qZKs3CtDDwqaxclWGhd1Tggk5bqX5LMkwSV/2elkMAkcAiB99
Ig0ivQtZLfHWUcPxbLIWXzqN1TlJweJUJ/tKW7wCz6FmFaJn0+3Gh1kmpu2Z/eZd
O7cdASIwq50blQhbIurzdVuIXSGTGeK7Jm6RuXnOec1Dom/lVVxzZy5WxOL0J9TV
Gtp632eF1tDtsEs8vw2qqR0CcYTAbMVs3W4Tl5JrWbvS5AydPow/Uf8YCahR2PFX
NamBNdLJBNcf+3TrXNYKNgt9ySnXdxypv9XoJWJOgYvRj9G0AvHoUXyI2/3OaChF
Cj8xDdwlOLVkn950xXc0yK1mGgluC6tT7NU4OpKGy90VPkAdjZgLOUf4aD/mXwjG
fRzzNDc/Wxu1fbSla1C/Vf8Am1iEEkky8/DKgiyX8GA/Yz4gEAXly2sDOGMNXRbt
E1aD46an1908BJPT2zSbpVstZQ2doxXerNPiMW311IwD9gc5iXPIwoDFUgjBS4RP
tnenjb1EiDZEL+aOJRBa6dqA8wfcb3bbRYduKxu5nvOLWoK2fHHl9mxCVTUmIAKY
7u8vCEbw8chu/tklVcTlN/lFDsVtiu/uj5l0MRg44oHvHXGd0gwdCo+gakMlPbvc
sW1H9fmX1aa+H+//9BObNx9158OQEc77RPNZkS8aGhlX/eVcRuR4FiRi9OyqvZu/
uodKqZv92LDP5eVlwpZsymH6gXDTWPH3C+/3+CLHomltu+ZbMGIf4hkF9ol2BPqV
QvwPsXRazcb1TYIzuEeiNKB6mfH0OTXTPox/QgA26cW4aewjt845wX21fRaT4QKa
l04iyK2BJLY+WaldYJlY/cdbDwnTKgXRMyxv7bJBboCdXczQj146VcaKnv0wHYuf
ER30mq0OictSJSR44CclAxqbZcuJ35A6QQGWSnF1icdcg8mXG/0W82QWFimTVHWr
BF2QNTbYBOf95dz9gXONur35y8dTwnjSOR3+sw/eebth/WaYPG10E+R0UOExILhk
MvEDoVFt+QIwiYrH9TArBTrnmiVWjWP6seEx5cYXDBEW/rFX7wm4YHB2HEfZKRNV
XsO6C1AULWEw3uCgl70IiWeJHVL9A+V4HsOvt1IQCfIDesbKSwi/TWQPavvuF8oy
Ar7nCWx+XgWIMssvjgJZ16aYTutO6MD97C4Ev+/3ytCWemHrOSVRDbnNJf5TdQDs
7qYh1DWTqyxYM83YxX6FzUz/dgSEO5DrznQQJN7UDeVTsfTRWE00w5m0xdvdZy1l
YIbazefHwlZ1bi8H1ZcZROkq0On0kkdx6vO26Z4izHkKt54KFXgh3ergs2sUePvA
IwQcZYvoAhSk3p0US3EEOsRZDjVdD5KyfAfjqwS9EojVNG1qtqM7PmAAkWdomSWy
PZPnZD8ap7NmANgYxOJiygvQOBOH8nqsT4hYpooqjetDlHq0I8jVMmQcqWsHXU40
jSpG4OHB6qFOHLrO/Ejkw4WZsWTOw6rkctnrIAo9FK13n3wZvO4/K/eSaLHfuyUz
NrLAWZ0Pl9Mko1ouJlAwkf2a7WwOjVr7i3dpiiVmbbFWxNBh8uqlvu3r3GDGzk9F
8xFVB5qWBlc+RbHknucaWilP4uRV440Nd1X1otbokli3BVhf7dARUryirwNWq9QQ
/Q0jkEBFkbdvayHekv8j8UmrIo8HtF2eJp1oDyNlOOjE2nt6SZDMBxssvlcHqqUW
hXa0nG/SS/cX4NXUvgfgazjhqUvZZmt5gdtuQrg54OiDjt1/WWdoguC2HvK9tmR9
9uel5RH8ayD+VcJH4ZcL9W2Fwg/foSpKDWKRrsuVMgv3sF3iNZ/KqZUbaNrNNwBD
+nPHg/9mx+L7o0vHws7Q1alaiEM6CHzeTw2pUGgozyUDEWonoPVC5JvMGl96WQ/6
M3uYvIU7OUAy/RyXspEzZOJon5O6M1yMYiVdCLQVqu3bGLoLtZsDUCudIElLTbzd
pLd2zJpdbHNC3kZLA934X74VLlKL3iL384EqVJRpW1UZvx7NQBdPJ1/yFy0SsSdX
pIECh7qQFe8GcP0Rlt2Z3jmsskJ6v1dlv9Q7fPllyfkn07RtrHrxarE+FJhl4+Sz
NNXtKS9ssDcVMcSAaE2vcz9V6xgVeoswVIku3dGfv4BwdqR3F4aOEx7ReY0usoV1
WI8M10bX3pALmHn7JJMAV9QXbfssCk/UT+Ajj9R2U6BhXLur4hsPea5KylMYo3F9
5zCIMe06noTRhnCuV6PO9E8ISta/iNxKVRMQvDABLw6BfRqph/vatBAay908vA8m
mCA3Ewz2NozRe7Me0BMcfeIyhexTdl9pHb+B1j7OreWgysjQSK0ObBdtZ4wX14Uj
CseAQNygGNeQ1CFBei0XoYWgsaAgQz2TuLUc7EHtieBY2qw5o+1gAR43otOZhW2m
8QB9//Zxpwtc1pkMwAUan4MEl7J/p5S+Sm+3mk3jfISJ8mOJmRVr0RUASB/FBpcD
HnU6A8Rjds60kfluySdw5QcQaQni1GRITWehm04cFyE5bh7v/1cI0vLQz/T1vwlG
9WBzxGNOb9/zkr4zo7Vy90VhaC+wcGk3FjvP/EolshjKBUgYsUlaMLYs+8yQsBKy
iXZtTpHRo2u6tdX54FumVPFMw6FLYBSWoOtxdnIoOoY/M0HRm8lZ4NV8Y2qsUIZC
mjgPStrG6qY3rLktIlpPHW4pBdqjxD5RRZxLTH7XflwlnNV0nDiK/qoPKJ5iQKEn
LGMTOXti/OusE4krYFrXFFCwg6+kWqoAT4UHpW+2YyG+BN+fQOfxq2cdq5k5Cozj
7KR4pRek+GL/ZVJhCA1kkMC60xDgn6FJY/cwSFBLfv4z4y1H6tFWXyabs56C2bze
I1O/DScVcnDFv34hRTdS2dlXpGWmMhv3mLoJlsW9XaOqF+1uS4G9Mzv29YeUT7di
s2/3YJxyNClCnaSKiv4e8bD23Fs2QgjgR3J0zokmBvc8LIC9O/dvLIdN6bEJPmtR
+1eMwYBy8Y6UioYsgPS7qGih8Nb/rILuIuLfd7QgfxmWyC9XDvxMS86LLLBMF57m
3g6fAtEWIuB2JQaySPZieJWetrKd/X3Xsvw5PACu/uQS618GezkbLgx3oASj2dMg
ZS12cjHuFvYdnUSnNOV0Qy+3WATLUCUL7w8dQR72/KnmnvtmHdq3zMyAGWLljUVw
PFxvO6Y7UfeoZEFmkqV6GesS4vX98Zloa9tP0+2BdHzY6oe9fowXk7afGJAMbEbn
ZCj9yxSp/X6mWQrGlJdQ2uy734tzyAzrIgoHvhp9nWR2qv9fhXy0i3t5cunafscI
rNPRsEb+gupG/9sCtnpUqbmMZRvARiYdNjWTHzmjgd487b2bJdgOZ3RC6VU0d2Tq
TzCdBCYeHzzm8Lgq5Vk5VQvTxEZbYu1xMfzR/Sne2BdhJM9xbRNS7DD6GHX6bsDZ
TteulhPx1SLhi4DYu3IRgRUfiat34x2+otXEnysRandx2N8v07oXn3RIOY6li76Y
x2dGWrGRl9cs3WnQSEumGW5LZigXpJTvvMO97gQCj3dukhsEkEJ7Q5CKK31fMZGE
0weYVObh7Zp4+dUk/2tMcC3Mwkp9ejiGgb0TQQYVZb5TblqavyXS+FS97KxWYyxr
/5uRP8pgawzbRMkEJJuMHSzVmKujVVgZQW1oBUk4oFhQW5fB6W/qTHzB8GJrD99P
4bKsgK0Votn7IOJzHbqXDFVW7gs3p8NFTB+SEk54BOzA+ZmH0Df6MX31dW3ifAwj
yx4U8DItg+Osb9jA5RifoWlxMuLdWpXQVhpdqeI6cpXSIeY5X3aOkvMt2/rvshEg
zOerqT9hRGFG80UVCw0BdIiZZJPh0c8pbdsuvRY2ZtFJz0Wbhd8070fRxZzkKXCV
BIvM9cOhkbo1JpDsg3y6oeY+4AVkBWQ7ObRsRQzY4/EUrJHQoDDLDUxKIIEBV/Nk
BvhzKRzCjlWKRpA5iRvycGgRLBFI1+GaJKyCFiN614ChLPYReqtanVeV+tCDXX5H
zPvrzxaQ2z4/a6zmsckjV4kHHd+ynH1Nuo+gmPIWojNQt/bImxpdZ/FAD+9XzBY9
gB0A26zlLEYFRKk6VEqDSmCSKbcSTv3nck4QQJdsvEGIzt/4Ye93cDKol3bWwuLP
ZC+mN/90nekuVkgooYeV1U4fTsozDcDqkIsP+0Ie3B62Zg4jQcE31c9bz15Ai/C+
FIBLOBAUZwAa+Sw60BQqcRImsLWkZEAwA5VilS9fcCLoQOife85fdlKb5qhdnWhe
4cl02TA4H3EouBeyGEY+WA5HWIou8HFxAo3107l9kNVBrUQq3bFPQhgI2Npq5X86
b84xDB5/Rcw4wgmDHgDNuVonf8gAA8YxVn2Jz27I3dMeOGxzFy7MycmlUOGlYps8
HxK7x0blcjbkB877Cm+hub+SPWId/zLQFM5GCmRmEJ61APnm9IuqTpXjxEM9gJUM
Pjd9GhaK5jzFC6MmQ1mMpTE3KeP5B2GBg7WikfZ8W5xfTx3OOOk5nKlU6Rvmxrpv
O2MR3GZlJkdVoASsRQXEXOxxOCLGG9Fii1NG54u1JV/xTxLoMQG0R0ThKSMS26GH
dkXFYgBYHQIXaVV4BpxwUDwbgEl2dKXf4Il7ceoUHjsWqeh7Xk6Gqv+Vegdm3Hho
oKgyVLxrGW1XD6AO7Jr1XOSzzWsQCIe6NTIqnaGZ6lbdxF584vUEqGQByvmU7GMD
rEehQmY7640MtGjZFsy4rpttrUsWlEaxrZ7bM7uvIYXAsjaCz+7hRoLGY/tj8NGz
k/qh16brh56OKGXtucFU/rQ8OUZ+8XSYe2TARvESLVXsHQ47BWXZgGfj4KlRIAvf
QcjA3DbXIiJYsz0a6qKBstH6oXs2dX3B93VMiocjkx9yZGzp96SOk7K9m4Qxvfcr
oJObeFI2NujGj6YWdUVZSlqpR2n3WUfBVbDglR6pE/O9JznM4UDxuyJALVPyw+uN
DibNUZSfKSxHG2lIRWSfKVLFEapUNKXNcnGQ6VyRy7Ranx05JjY/B7lL3YyZPUcT
vsKPW0jHGZB09NrEZR9G7AZjI9btd/eQtCreJ+WlK0gdv9rxb/7NOXpa0MfIwEJm
JebpOpCkC2WoT3yp0sTnj0PpD2sjDipi9JhECPkOARXr+xSkMkKfReydkW83ApOk
sNBsvv6QItGl67S0D7GnCedGIT7hdjyZIiBfKxlryNjk7BIYtL41Vbjrxpjh0jaR
v8g+hf1ysQR5AS+nY8n02Rh/AuJ4Vr1VfbrF23ml918ee/tGK1BmgU8317W4BW9C
EM/FyqoqN+1+vLjcO+fKrK53caYcB9rqrgzaMCQakaFQKjW0reKsr3rnlIQEVsLt
Fb+Mt9w4Me4xNTokyxN5SPedhhtJDH0chiKznVBYkmrl9T79nspcXsFYs7S7j+jn
cpfMdn06qS9gqdx0r0OUDR0lIcGd+MCJuaOCquzJtVYo4gMTLluXwetFhvkT7v3Y
meHvjghd2cspE8AttaPhz7eOtoa4rguqI+pUQB5lZNcpVPlVKJAGpFM54Y/DzmVU
yyphJWty+04yGDbSBW9jdf40yYVfVVp2DgJXTRy93ZBKM4n0h34E2p7amMulBkS/
QQRVz6soyQZwH2/AfqcmDyyH2FkfiHrBaLycBcR6D1EoglpSmmYDMSs3K7OXNADo
4Puha5AhtykUo0fOcdbMWjq+K7qHctoQHN1opHkKCgEh3fLt5cWFo1zW46zRqjyC
UwCb3sIrmb59Vgpep3ZrFtU5eV+FTJdeCKEivT1Rih7JUFewMp4CyyegqdYHbklk
lYkGCMVk1X2cIVomVhPSyDOPktnSU8PqPrmBgIuLLnEm67DcUVPDZpXW9+T0Ndmy
0l00bRSgWKpTNJqU9EhMWMgOSICAZG1zH+uA+ZQ4BXmtuUPnK6NNsyBABML7IkEv
TuORKODXcPfKCu9Ad7dhudTDZSNFQTBx7pFA9YTqoBNfkQxOr7TicE3q8i9C2cP2
NUgEi9IjJYIYX98mH6lyUymkxXfvsqa5oGYmkYdtcDtxswhXI34dUBMa1z5LDLtV
pNPmBknaTqEUieQra96dyljPAYkXck0Z3+MyEhyacsfjAY2jO7PKPb/v4NNDai2p
b3KN/APeORg2yHwf3IpciNA7OIIiMPgvlnKrwd//Sx07CfX0+L/dxTIhrDr4YXdg
Kr9Vd1v7HnSbmZTBL31J4/XLBNRD4h0nus4WBI4L6En8S6gFCVhwYxZCNiRo3gR2
dc9dGTBE/DbSl2mHesLNO9pcxCtRPguIZqKtpQYzsBrLP4gMunJQ6GHSE2HmGT9i
WtUmxT6aOtbrtQB4NpBOcr3z/0iqZlCnWysyOMdICKCvT4ZSE5rD/V4m8V7uO0td
eSlZ3setmS1GqD2kiooOGkKoPhsvKiaq12oPpNYgVYfNcDP5NGZqjxjHL315c1xk
N93JYjsNUTCDJdiwevoNQ6Yw4XlX8gB68rI9CEC5ZoxVBFDMckugECJ59t0l779p
u6otXmaZ0f0FihtuD9kqwCaIvI1hCjHIjvIO4eLR0eqO8hCo5SK4KeM2QaIV3fNI
zfZb/Skasu+sdXEoo3etvuTkeeWt+CCDxzFuuFKKdb/Bg36MuDc9re2wtsgHCSu7
9GHn0NLEPB3yHCOexw4v5fiYMToKX/qffA6nQmqOB/o4mh2ForXuE7v31K6C9R+P
CfOcQtym6FwSyHyd/i+3eHkeNiiiURxZjPvHBgUFnPkTVlZurMT75lHofZQlIjZX
dj5d0qHo3cE3VUx8yB+dx1vMNxpW3ozEVIce0XOvoA92EfMJkdktcvBroFaecpIV
8PsynVdJ8QFckb1olypOlEeyHa3m/weR68heiHNHkd7f58nDBPK2OW7QnRuzI5HP
BbWosr5TMomQLrI9zVyorrQaqg5h4xo12jS2+WF8uAWxRzgP3RX681umFsi27WrS
vWl6LhUp00n6YysQ9lnahfa2NUjYtjYJyaFk+jPuaUs7Yt7FIRuSv8Hs+5hvZG6L
WXevyxqgs/5Ex/P5QArB0Dy5HSaltdcEflUdSqkHN2Ti8KNM6jBJ0eKqe7RuQVgd
8yFNv6PEnvuEeWxiOIk4JDlghv2tLt73jRVHvPRErEL5OW1LrLWuGFen+ebO6WP5
b2kLTaDyrDuh/KIY/EmDf8MX4LYMyA/yoXJlPHc/+tmBw7DNn7Mh5sOCU7RT6zIh
ZRJAz39gmZeD5muVHGIN/1bsg44pKgAvrw5uz/kQ6LKtDK/+i5FnHLnmIHIYwWfa
K/nNzWDgIqnqMyDVkYXSAzZ01Z5cQxAqVnErjEvEe1YtScZi5iE/a8zsDNjLBzdW
iizhR5l4G4U/Jjo6wOrJDuF4tFhm5MZSmlNQP4S5M54DTb/S4/qFil4A+s4xZCj8
dTkOPkeIcEHSgzLavolyQD8hxxAgg0Fy05auUzli0tfaQrgfHvTjq06RpjYroJFP
WiVx+tnRaDO5vXnziWdiCC13QFuze5MkzfwHehFCp2ox9aHdsr9YMAbL5anC4v72
3pA9Q2qbUdJsxFaRvzCWSho3OmKUb5CBkRKCgZN74tFVXEtqecz6iEQSJZEqMy84
bUCTbDvnELTr3prYXQcVYh/d0HMGbjsfRqrYk5RomfBTe0OuWYIZGhDCXzO1fD1G
P30bknF6Z1rrNHJ66oPiUI8qxDhd949mHizOfQ4+cJx3l1FumFc1qlrMpgM84cjv
cmFtYslHXWA4/o6s5miv0VjwyR7YgfqWs/zslRtbNrQ9350aRlRId9qG2DZM7xbk
D4tc5OsT9cCIf3KbJ+jj4/IAXQfly0x5XyOm0h3TR7HRnMrA51AHjFRxRdOIYldz
NqHTSeiusOJVuiDL1MV/yP0qwSQcEdut3np1yr0bhVVVbvXiwurE12UIWyS5mIlU
OlQa1pgEIFEvH72lDQkdV/GlLSvCKaB5C0cfEWsey95/cYB6qRyZ5MnWIWhe3ub6
9Q22oYjZgzbf6JHarygKzi4Fr5fGyziZ+bhgbfSxrLfDH37fJ7fH/0oG4lZEhyBI
CF9XBRGr7JCh2OctrW3XhM1O5cB5rCjUCABmYq0oVccdHxYxqNIyL8ZA2jlaRWfd
yeyH+ocwidznrSrSsRDRNBVYhMFdtFKECtWsxo6ZodoNeq7BpnhapY6a6FVcT0Lf
pC9MpTKJ/iJqyLW6M9J5pqKBRTaq+qbSDx0OSvM9SXPqTbQfizlPZ/DIBUrxjlfW
l/w4bReW8o/MCA9K0d9R1BwFrGc6kVTZuqjMF9VtPGYqd3HCQdXI5NHoNpMQ2VI9
CVoBDV++kvcbUwuHi0UUQfqyxOSj4lAWVAfCy7ghD5odKORSQ7/S1yrrUygFTJh3
y6WYNLlFGLfQYv6Ho9TdUyR0QtAqfH7UA9++LbcEm0s7dB9mUqOTLCj64Uk8VamQ
dsNmKBzoQxaWjr3uAwfX6zsjHvJLMJ+2l99do31jC9lF9WU9gr6KdHZg5K6qMUxs
yPgFIJPDxDhn8HgLqrgdunneyIQmbrl4DMwES4cBPzxZJbbnQVelryWFzUJyvxLx
flXKKLJRkOLYPdUUfu2LKHtNa6kDeNcV9emdroNeLJw7qECd/C419OtC9ey03MAi
vx+eX+xsgtLGxmEBBHH8Dtv+RGlx/57s7ZYcSsRFkjv7leVcOuN0dtGaYFOn0otI
bEI3SEg4yJ+Hou4d4ASf0smT43a8OULG82Mm4yulltxbkPvjrOKnW8dFUBfmtPwf
ZR6szmzeYVdjfxhavyJ4nU/uGJ7bth7ZS9GvZUdTHxuG42EKsGXULOu1Byo+0o3Z
dDbPCzcCJL9sS1akOCGNEwn9VYYAG6x0IPHoYZUfL3Y4btl096FF4NxYtNi1MWIV
l5HLT8M0b6+z4UGW0ClRGveJEHEJTolhImFk2jnpsKLDSDY2AD8q/4UBBqgRPi0m
v6qGpHfPKqQWvDbTtFBUtGoNZAU5ZsFayfH0t2YdaMkgbMLVAqYByhEuebwrs4jI
o71bfvUUhWc2eY4guFsUgfq6SdQxiVlXWlTaxqQ/W0hIO5tK5rWR80QWM6RyQelf
PhA8ZPgV5sE5g1oVgOy1AuA6mFqywniwbT5trVaaX51gWQsV+UDSlMflWZAj4gYx
kU5ICLv1JleDtlTg7NKai4ELHepwVQl4MqWPga2Qo3B12w2/wBCO7v4gwvWY1Q4D
vRxN0PvEmUfMqrDMKjD0loiRkaNtB0tHRBKFP5C0CZDCEQVXp8k7Rs179+q0glYG
q61oIvJzlNej4FMO4THABNjeGJ+yNXaILSKz+NuR9ZOaLUBfPmihtrIJ4QbjsMkN
PU7WWRR7ErTCpZER4ZRozcL2bjfQUMlQQS/zRnYhH48XNaUXHHLbXXdvUZF/wUkn
enjKb4StLMGRsClCYKBW+au7wIXNlQdQkK72BslbIrsDYnW3s+8/L0901rT+RuGw
Zfysf1GFjG6mATMyMBaNpalC23J4Y8j5n9Ssb3xwZDP4TI48ifDWrat+mCtq0eKM
lCE15zK+1KXTYoJzlw2UsTcOEmG0Jil0Khy712QwfzE9rPmqlLKpD6zetQXFSUyA
K6TwMCrl2/XDfLrIoW9gfserlOs3ndJOylU4vYCdZ+DpY93d9W22RYBt7nc3hbuG
Yjh472VIWFN4rZNXlJagEAAJ/ZoSfi19EuCsjKnmSmHu5G36xPnM9ZANB0A5TAwx
aor58csXdqKxOuH4RjSLSukyGKLH706wSRqPz5a8Tgqk+lmEhhSh548x0IfyPOfp
hMBuAO5nw6THlCD2WSwiWjn2zd/HQyagphExqCXqQL096vQBOtiyMdncx4fGM7wQ
IpmP0TGvqPyLzYR/Rf3CJOqYYF1BVtUntypCDtRa2A0OwqBht42OF4cFCVvjZ4tJ
PAcPbjl2QLJJr6Jr+eDCKIemqEced4PUcjVl1TX/ngD3fwaTtkuLlAnfsXx4CUH6
GQD6Bqj6QHCt/LqKVqgftolQVHREpXIkbmz2qyjF6FCJM1vxCsbxpceNPdsYNaBZ
rgxLGCKSjEWRULApo+ya+ml0I4s4zZHupltLhDh0uJx0GrCdKXKPe/nZULGkvarR
FzvSYWjRAW9ZGlPPwbjWEtgxCcW3yvaIV8E93E6ZO5JfsBGMG5PysGQ1b+gBmQFu
kbPj5H1E2C20dQgh4jtHLm15IOXdzIlfms0TnFpmv9hYF38r28L0/OFjAGx0Fmm1
+iWVEzcHS9iB9O4Z+UMNRGm6MUylrFARAGxoeupn5Rs4ygzciMR/4kafoeoJnp0Y
bzivskjwcGjZysipJFMKowK7OmnZUkD/SblVOaqQ3aWzlYOYYN/HKzAeOM1H7e2R
EXW14pQEUmNKfwKcigYYU69gkJp4l+HJ/UvoEXjdU425MxhNdsTO604Y9Rr9+v9v
LT+js6l9V9bQUhXv7G299Vd80zJBEBvHpVXmtqMrSvoWmu2oNNOsgv+rgImuKToF
v/DzAgU7dvU9qUH521YTXQPY68Kp+6iIqTOELa6Y3/IAjQ8Qx+EQ9n0k4YtASz+L
NXp8I+N3mCJDpRUsn2ifdAoQB8VCb21zWdTqo1FYAf3uLrC8AG4Xm03T43Jv5kS2
EgkMPhonsKLomlGAUvQgF4oNywWJCfXXvCXkUPP9AN7nEQrurK45K7yvV5TryzhX
EOPcTlnwbJY9QRyBcp9IBVR8tu96S7kzIUp3LbFvzV3To/Jsk3WsQSIYl2yLQsR1
sNSLCC0MVS+WoXOL1z0+BeJBu9ryAOKHfByATe1/+c7RX9DZuI3X9JqXJRc7h5mw
hC1e3N6IbyzXl0QBr3KaWIzgF0yWMBOsgnybjwXutMG12aC1+LfkxuSIaqDKQrPd
7LJle+i6YeiByCScq8DPS2XazL8+m8lnASkRy6GoxaQG4tuJuujSJcXr9yJwhtUA
yR0KDmtqAVGcjVSDD/D1cSfOWBiwgje7WIPAgBM6AUsf2ndfLMwIr0tY7c2ULs6X
bDx1oKt3FguENHWi6UPArVPJC3XhQSA6joan2rdpntMW/4rBrdfOHQG6Br7TDdbB
Scl6BbPXTFbahCInoVxca+flTQ0PLuH18SiDk4pCd/dwphwqlrdNyb/r5iu3cOa2
7w5lozZv4Cm4tAprMjbKjU6JrH1knpV2D8HMcfnzCryEbHDpBE8BkdZ2UEfN4rMO
el9cXgEdwlE86ZiNFs62B3FLMkGv4irNj1Eq57X5p5VFZ+5AKKDrNN6yzkzZS8BU
d8ZHFcQE0hWF4nlFZSEqFVOBdJLOtuuj0cCqpwOO47XZpaQnkuVtolYSa1HYKovU
E2vhhkHtgRwZd5h5EJqbL+V/d4i42FfkkPnf9FwmJ8W6Dqbe90KEQ8lKopyUFyo7
gXd2pIoBFrs+xFwDcFoG13TjoUqkrzbb1vpxu3pBi9YbxvV8eG3QJvTRyOmgBYzu
+saIxcUHP4C8GeKEjKzwU/+wTK+j0m9IeSk1NY6+OBDOL/Dm9iToWbJWkgxP9Ofo
nEY6axNv7PV1tuv/scOya4VxBNpP40ZYNYK6Tk38fZKy0nRrO5rW050MSwr6nkk5
wd3wJ8yqoZq3YQmW3+RcCToCDTe/XHZl2l+eVipuz2ql5dxiGAG1hpjPhsqqp4l2
jfUc1Y/xIiJ/cphICiJaGDSsAT3GbtLzBG97Kg5CLtrk7nX2WrWT7PJb02yNlkrh
u4CM+vtl43XVCHqD924v+D23nCjjw2T5AnMb2BIkKOMnP20lJMPRi89D9gMDCY7t
JcLzLftCSxS0dykoaWdzenI1g3xkzQprC19XzBHr5/Yh9u4SrolFOgYvknX0sSYv
dW8Y/KxYD0u2CiqIiFHeAaZc+OVtyykxhnG8X5K6lUuS7v6QmBLk5AbVNEJ3yFsL
8VT9+3+kuq6zZwrR/i2vtaDZ8LzgE0nCQBCrUZiCt6HGWwSGZ5I60OFhLlOr2Ys2
vxSNM4LFRbJf9tWhJg7+7RIzx66HBAtWc1TUYgyPM3g95Py2iHekPV70zQZxPfO7
wuLTD3Cybo8t1SDjqBYiHewp4BWniy3TysvaiaIzZJbNmXyxnw1FcmU4vFlnnG6V
7lWML/ASn/rZl3hV7XvnucV+oP1wa+KU91ei8/qQrveSL2P7hugJKDjxKnOzsDuN
yCCUzz1imjtLzwPkrPuehmnuF8EbLVhR+C2ALeUguDehsd81rKsXOHNtHCT3nCIo
nLbQjGKgTNq/fxfKinsRlaTDtQ77af0mCszwu+XBHh6X6Nlf8LsPZ7DxX09WUsSn
qWlVkmDJ6whs0VBmPNBOISFhGczpfCA5zBhUblk8z4Qx73l0EN7HROjeLGtjogzd
WAllT4mjknODHV+FYJlR8OiYSRYaVTwdbDyMZHg2gxfCxuB87LVIxPpYirif+r9C
yE+Qf2vlOmwVxqurpAkIWAQv6+lOrTj+PXRW8uV6YSaqg4AzIL/Lso++i84j7fAR
h9u93HGPj7ZKKhGy83b/s8RzBOwhBvbz1kgcE9vBILchWYtnXPPbIQd/WeRlqwNI
HXDCf0a7W7Dp/GGXu3vh+C+4rjGUUZOwZS2qMnOUNHSiIHClA9MReA/3Z/LRELg/
FutoN9Qeg57oQKG3104B+mCTotZrbufHLPRDaqGlm6smiGgIEVD4GvSega4A+69+
Hnt9/tQdmzWYjGfCwre8sJ6xm3LdWPkO5OyfpsVIf+KkDDqM4yMpWCBuA/+8UFW7
8FnGFjG7YIhNcH1AzucArAVrrLHZwi2gXZpcRLJLkLDg/6Vkb/NY6AdtR0K/DK1s
RwAG98ObbF4uF4SnLCr9yMOiBBoZeMyzkMixLUNe2Tq9LQGf3Hs5zPtuJmgHiv30
NXJ7qFsOOv1woCtqY7urbwKAa60rRPfoPZhTRv9KsvmPHDVohPJRJ9lxoll/eyfq
7gIVYZrnh1H6q/bLn+ARMZDBM8FbIshCdXe87qCQyRIUlhgZC7qWU2vh7jl0sCDT
ZYD4lyR4AkmQMQSMvOKFmCWt1oTo3GWL3VSxRG9SIjn1cdh7Vdd2E7zv5XCM1sp7
2ubIrceiuacblLNY4BdeKc9n/EPMdJbyNsjB0o1aEX2uA7CsrlFCtIrQ58jZfiBu
D9qVpamaP0jXg3teICSknZExcelT1xXzdl5ENYIaAvtrdbePF9C6B+T5iiNXsck8
zq1zwcVMZkWbQsVFqkzN9P8q6eUawv/qJR23lD2GO8s+jA00AwBsZoSdRInKYpwG
kmnGDAfNh5KTZSxd92T+kLrGjhsIWfTxxshsa1yPvUGfMylIrM65/bEtpWay+1UU
86GdejrhklX+c4sQgCtadJ60HtYuFE1Rd8KtuPvprMAQtHnzDJJmgN7uIsxBFSUf
pocE1uPXKKRmbzJNSa5CSVoY8chsGxgHywvM0BkVXym98FiTvGrRq0V9pDCfp4yo
ok22hIUPJ/yjSSziGYVCqUkPitq3nJsJrIEkUFHQPxv58PvHpOliXnVzeRRRHsKc
mFCZO8QfnfsSs7wytJYzsWsajDrJHLUjuZlXI8vJ0yToLXSCo5I/8IHYvWarwt+T
J8oXq/kjDpG2SSwCfw5atPImOO1zmkbCUEBw8xSVqsZ4S5C9R1BBsc9kKjXGrK0Q
f66i796+wnPT6Sd5AlK1CNHLh56TyTl4IfYzXDDVfkZKGM/LeL7iWYRBB9Qt72GT
MVWBEeAvoNbLkHKUXJneFkeKQg/aKKjTXTM9Ijh+jNEDv19W3zGxbdEnuLWbtv7+
cUjdHTBQBIca5MikEA1lv7qLFz6J8G0kBKRniADvZPZgr6gAN4pOXFlwxZqK0OYL
DgCtTiD5gUUuVcEeol45j7+Gr/fBy/xz529Bcqueoh5dS9YmlpzV0QlAPjzd9yTY
2CuPESOGTpBggyXWeSmNU9A+Jju5vrTxFfqNCFYqAsoVTE+qaEPawRLDJMd6apFT
I/gQE8fo1Kg+cz1JuvMRqXvD4yaDfp0COpEQaPLFX2THoJSFi1qhbCEq2dQXu/hy
QX0Em52cS10M7Zqv89LY0/kBgFRej71mKNrs/XfVB93Np1MFtCHxBHbC6kRdeuoC
HAUf4wtVzzRRXNXbL1XIUKy6Ty9uNj3GFM+LCMRa3Z9A/2FGXhUdJqps7/PpmV+W
k0efNCfPQJOTzWh/aqubVCH3rofsfYsg3Vi1DVZ6UKCIcWIo/e8udRVnWHoem+Wt
6l2rpz2FqHGuToyDBXTdwefnb8hqgi933fn1dXbUsvw3wce2UGynChLzhIsrdwx+
eRFWEd0N2R4/Z4FL1rwO3eJjoiCt50v0CSK+QdcLyGBeaKDHdjqR6QU3P+Cjka9K
BviHiUSMudso1TbhqK+k4WtOVhJ4WX09P+vB/qnhHflmPi75kv65AJ3m48rDs+VE
glZHJcgGXinMX3Va7jdNuNNkNLyj6LAFkrw27Czh8qevT+cLipGvt377DU3h0T6R
QHTZlqxKd0yk5cRImKTuDb5KeygQtcxQQle3QFyMlngudiwKQcB5JAHwFeF7QHGM
KmjqO3lhP3S59TxOmVyFHAZzCVwl7adikD4wZCKMdhBMlOIlcXByMRI3Cu7Yp9ee
EKLArum8F9VbYoIZLvb3Q3o4kymZoJzRv5Hd4iHDMBv7sS/DH2ngz0z+lX9vncBO
rob5fpEtKYJ7d7uKqMjS1lMOwC2BICmlrVEHSrVWjEUp9BmpivdTYGPp7Gg1dnme
0N2F7THlV3FptJTeuRan5XwadIMGA3EslHqWgyWI7vBXnedwl7HwncUFlo/+Fyrw
BYX3kh8q0HYiEr/xOILoBzoFKQO9A9KyoswIWwkFwjUnG6ZYBvzBx3t4CwRXzZHG
YzXDcHwQbggcQFbKcPkwPr5gmTpCkLDN5KPxj0EzORBGzMpQnP4/AK5uQzxQRwCW
qr3zEXSEFKktIZ9qTnIWVwdOMOw/MMueuXOa10kEX3YqbDHwCJ6GSyWeSuaFCHHP
Tj0g2r9VZBoe3Gb0gPomHvhDrhVxOKoM3r/yw2HCVxlJ2aP2kXGOActG3FTUF7F/
a87Nelg9TBKM0qatm1q9mBYvNqxUmXrDooOuEV59TVFz6KwvOop2iIz0GlSLg34D
ZjcmujdM4QSD+xsL0x9+ZZ67KbLDz3D8LlyQ8QkRuRX0PAfkGVV/ubGxfxP+lvq3
TvoXPZFFDimUF8J9KtMzcVC5X1P4sMKEDfLtguE3QqV+q1E/Y1fY5apINIelIRcL
8ItRzUhieUoWASpz8l50JOMpZQk0vF+olpOsTn4dS9uuDmnQ6/OA6ytPi6BiqeZj
KyFlBXeS88kHZ8ESI9L0/g9+xLrDboVlax08mrQS/xd/B7Mjzp71Kt2M2tLbBX2e
LrSayexrVea523d9CDmn6hHLhKrd2msLqdPvXofYvRa3E2Y/QCMBsmxx9BEJkE0p
VcP/fnWmmJbLU2QHQ0tzH3UghxfszlDw7MN2NaXxbtaFVBPetNnbm+LBtaPaepkQ
nvRTC/QLboohZ9NhfqeS6GQKKEqLlCrC7Gc2x3xWNP3KaRrOVUmJxwuLdgRDTAcZ
BPCIeV+D4BwMo2ZkdD47caDNn0edSDSk8aGr/x7ji5AhfpmUPdZ7848Biv7Cr3d9
Isi6wRXaLW/bNIrWgfHigSAJDLMIuHr8ChwJq66kdFZ64ZF4AD+0oWXRSxlmPG8o
F+07gIBSO7jsjlycI7jSvgJyT5JVrA1OxmX2FCa9InPJ9b++UzF4PNZkT1wVAaNV
E8EH2qeEhz/Zsg3l6utgMoE80sU9YEXgB5p2L0mJlsSQULlNGIYn0jFPPd079aTJ
XvSdvzL/XGmJQoNIdurhlnzQzlDojx2VeXiyGvw+Jls+7CsQn5v+nIAB3LGuqJbi
LDyRFRLcjpF7P2GTFbudcu1GZwhRqHMn14m9bR8isRVngQmo02PIpTViN13qDKoK
2guoNicUUOHtLXa5zCPeqa8benecKofjCp2nnXysE8ypUuSGpQ5P+BxiZky/yPiS
XmBMEf9xdJibtV46E8VfLzfIqrOCGK0Yoq9xWafEnqH3/z/dU1S+BKGp2PCyOAmj
bShzGVChz9lxPWfCTIekf0rG2VbfIJLqH2Pgti1Qq8NieTjIMPq+sH5SjmFaH0Gz
n5LksmUiJ1+f7EXFtn8xN2j9uU1ACHuEk0ayYGEXHcGup9gUB7WoxDNI/Tl4/SSe
sf1ADeIaGbuZbhyyW0RymK1ukslyJywUCcNwtl8A9ofalkK2UykG+xUSy3h+JuJi
DceTVNP6h2SVBhiYmVq8db8RNy2J7rQY1CCJoxyXCh4XDewlhjJzgPdTOzkMndK9
m8t1ADxexAxaIz4e2bJk5YINB/ed1cbmgSvpAOBtuNSAweUPZaEgItLP9k1K15qo
n2MhIJvCLd3jw+G8MS1lsaPgz2pUJ4EGEmySmV7WNKbFRW2s1Qdw9HroW23ca5Wx
WXRy5ax4P9ui5joBBSJpXBxGFX6BireiSKey5SEgtZFcx4H9j5XdiahRIJTOvCXn
NSZRdwIIjkXAQ7IJyFG7JjuoI6BZUEWU2XsK3nP8rhDAGGLo6vgoCY/CQKLH9+3x
rHQh6IkdFCWB5k5guajSGzQwKGekReIb+4xHuRg4MHQ5RDAFw41O4Bw+gDF6OTX9
AQi1al8GoK+XCCvcz6Floge2EYY3uWfRvJKA4Is2DBcVARlsZzQsq1uX9NMsPXKJ
CjCAgygjsLPMq3CgrQx6F1/xyCwYZUgWWx/zAXV7OAAuHtOpbVymMXE+UsqQAfcH
dcKXgsBUm82ljbPSnzInkcqqkZK6yCqo9SrN4tA5ClkmRl+2l8BF19LbVxPaoDAC
zAdPwBeWnMZ0m1UbV+OyEZE6FAuIiWizdAg11+X0CE+erZu+tzzS0V0vILwFBxLT
rbQASglNV6V6fwQR37kERzNiEo3CjZy+YBU0ozfcDsoAmBNnOMj6g4MEfDpW+L7k
qPFsJB65LZyu76giyezPjtnaEKII7M8/YqZNTFmW2gNgzTKWrO/GJ/Xb4Poeo+kY
p4mA7Gsr9USzDGjzJR9pL/OaXoJBHVy7o8pm8NOgrNwmxnJvPqf/rYSY5rkJbqxb
EMAWITiTvl8aTlGhuet4gyyer0Y/2CaiEwc5UAfxc102/FyAhZZ6XFOhoU6q3Miz
/cGhFBku5ElJvYyg2p6OV/H0TQjoGnhUEaVTAEODWpgAoVVE3w5++Conwtjif3SY
IwrZTd1Bk21+qv+XEnaJSzFX46+D+AiX4Jd/lgmgfVlLmtLzA4wVWdgtvjHh3TzC
wLovAx7nHvtg+SplTKi4RRAzhYXeYmF+SQC3YwmlrZxTeNcqcrMfMrUvb8XW8oUI
bLdeOQw0DD5ORx/rwHE+CWnGNvX9NgsFly/aMNrc57u5gcUCGeoEVPlR+ONAkCpt
YqunLzN7W3Ge9Jha+zqWYhIzNnvzg2SQS8Kj8J1PNQAmjOmKZob3dHlEFb6cW/ZA
0Wim4KGl63BVtcNecz7tUHFAvlG1EVX24RYxtiq+6OoWTIWIw8if8IhiU8raBfrI
aSFAdFAUkN56q3bGPbaRvshOGHb2wMHdLVQBXsI80WCfm6FSVsSxoYWBn7dUzbLc
QJTXKVOsm3dr07qh+GvzWKgfZXxdKsA+2hLw8h/SKCzUWW55+q8sDXm8fTlf+w2Q
KklZxy8Omstlvt+DoUEqIusGeV9lpkb9b/LSwXWMf29Q4tCEnigtb58nuIN65jus
JroEZA6ib8l3TwV/RnVTFf+KusHjC46bwdAFxPrISwQ1gojK7bebkOXyXTxhvSit
CskzK+8kPIH4W99aKN5wUpMrSZwmJgCNFqCRvrCLfGCtpxyA9snRCBmvptS4bjjX
MQ3YvwdkJa+tVDFJAs7RYHg2mff1w1mdNjpGfMZqBU1okdi8BEVJh2iiXdSMEGpn
FoM8V6KG7xgnM6VXsxsg7vL9dra97IxhOQMlun0VpmSs3K8RPbvNGyGzLr7tsLrs
3aQcToLoU58ZqIoO7ydUA0pddF8zGMWuHPO2JmkSB8gId8Cv+PPnziwkNC9cE9Fd
8clvoQA3ptBKTGb62uALU3gsA4UlDMcvEd9bpEnqQ67YpuZ/0eWv+lpRSUDJ/kHb
clSDgRbGQ2z+s9HgkS4i5meFNreunA9rLQ9cu4QXJ0C3JVn2TctptZYm6cCQ9lZB
+SrtZqvLveYQzkqClME6gArvcPOooFwoMmZtA7L0tIT2r9iYhNayLpnIUuSeaN32
2NZ8tBRH4X7KtC5zEPVL1A7hIVrOFhZS2E6bxZ+P+axDT76NAqta/RFTkNOXRBmv
cVTunEEHfK5dr/IuTCH9gwRLOaNVMdSNR+jKFV2jPNs1n2gw9RjzuJjzwVbiE2Yc
1iKJXnMbMegBFaS7DNuTs6Ms9Ocjy0WlfbnOLDqqhm3m/fC6Fak34KSqU2Il8RTQ
07RQ+wqZ5XYYACQq39LWkHTmhngwzQ1BBvgFemL731cXWKYroIC/8622q8ChHx+I
l3Pu4Wvkywp9TlhbsjnWINql1VTIpcWa7caFX76L2iiLtSEjhUjRd25tQUqQ2lOe
W/1gSHF2toqRT0MwUtGNdzFbecuKtXPNcZFvXMTuKI6Nqp5DKpCju691ymuoZlWA
Byaww3l8UPBHY4+5uSW7qgHaUsOI1Lr8dzQcRQ3gRpo2IadBJRTZ9Rf9LA3xTAn4
QY4G2OEyIJKpM0RvP7HLbA827Sm4iJFIEFdPHj9lEaEhqGPrungDHTs8qsgXDa41
JfPZMRF+zYg2loZhFvgedaXFWyOIA1cCT/ajanuVFBfPHilLWYSMAyCvtKDBPYOT
bmS5A+xhK4Zf+wqb9UnDOdp4d2TNpElI5yMRQz+/je7uJMJkVjVGfxvpWvkdWaKJ
/nfIx1bIa3olk9Mmdeg01sUJUY3RsYoBTIdOsRZfNfHIKZqyAJfFlO6fcQA3A6Dh
SPKyG/hhkcHYi42S/IdY4PAJa/dm0u+KjbvSI4Secyvh72VZjhgzmKycT78+Y9XQ
6sl9T0XwR37yq9ngA/NI6/P72xafWFK4HvJeHWqwuERkM2amRffZcOMaNYINBIoX
kZxD3OYswKvlBIq0YbWc71BXQPGs0nPp5VghQFriIJVVBCrbOfSvmJlvzuxyvloB
W4YcyfNAXmcV/s56mYvTY+qX7uzthDCna907a303cVdBSShudU4KzrtyPGB0jCfh
n+SlotTY81R/GZcOQQ8wbOnQZnFNAI1Hb9wM7m8pGREUq16P7eQWeyBMjcqbbfIJ
9dxGzX21he2kBtiNp/u+Th0p9LFIi/r+dVFJqs8l7rPNzm8u+pKBYTYlzNsM9gwh
HBi+IsnhSH/MNkeAOLpA+jr/y1oJeESUNgew97YrxNxfxMPGieCZNy5ZmdTRliYy
YLL+xSplcV3yExrKp65zb/PKMAG5uDu+gIzwQgD+mwCkIKnRNR+crI67VAaRFZ2/
Str+61F1J0ZDXRNNNTODmIhC96J823Yzl52FQCr7Zu+OY+99jKgLM32pYvIAyeXk
dxgek1AijZIDxjaOEU7jGt3fQvdBDwZAZqzUlhmpG00/W+ll3MpeAC5dg9RV6/Pj
NS6qF4bIxuKiWYfFiZEZZ8XZxr/VQv7JOPRdl+bSz+SRstaP8sa9/th3INyoK64F
RPtKScXSj3b0e/feQ7MmbnHuL2mxtqOQABK5hDJHJf2kXGlmpoY6BvrAVbcY1oUq
NaaWHtXYdvLVtPbpwrTXLe5HrAdKhRtlQSWXT0592bPCk/s+kJuhjgDSesQNM4GY
T0moKRr7G0LwRCW2K32CqwAkKmH56RKUHxpG687fGdcEqF5HASwJ6u11+St7Ct8H
gV/2rRBaPA8vmKABtrLG2qkio/FTgvEgbXnfBqzfn5kbnhAVj/SoGNY4/QM2HscP
r5kuebg7yoOzTajUPxtE6aV5atrIdmOH9mqDrK/SoFxC6OZghcqvSYmAFrLZCRgf
FQBHDEq0kkpt/WMeokBKcvoEESPFP7tyRE0DiI7OJ0InKOGi+WsKfugJOCg+AJ7N
O5qraXkRnaRXMERZ01sGK+AvgN0mB+lEX0zsFYqmCe8Set5x3Gz4lJNf4soY3hpF
fICK5GYGRk/wLo89XxCdtwhHgttsNUKKQak7ToVPAboPX9g2x1tqm6QYmpFuZjFe
8smgxxbHA0mA92O7xrGZ9FGGq42ETujGmfOmcYx1d7cLTVMWM4TDa2nxWIp+xd6Z
659PEuX5wpkd17VbA73UbyQoNB0LLK3oqK/G0P6x9LBejuf2PiLftoZUyxOXWmLW
9V/eFBPn0mZweQT7fqHgroMgFrxREsxOXDaiD0kj4364SE9ScT7jfHQKYOLC5ec7
lZQk5viIcoMLgV32PaBRkJMsptsKF2jAz6e0s8Y0JTPygWJY7i35HXoP2b9NdWJK
au2/Q3NGJEnV6pMXWP/LtLhMsWGRU/OxMKWmQJKieYaKEjP6wOOZ45je1Vc49kdQ
xHHyPBw7TjoSvfatWA9p3rtASAFEVMkO/tn4/TmufQJEkQ5A489mKqMdIsKf7t1J
j7odbd29Pe2+ijDcYqQJSEVeFRqtWKJftlT0CkXlBLvGiVNL9chjOO4FPAs8nDo7
7XQcAVl+JAz0YIRJECgNGTPWvnIz0eMekEOj171gQ4nb6L9H4Ywv64hBSXps3Bf7
sWBr0lufUsJFeSbR0NGl9dsXtYeYffKLLY0iNAJyPURiEM4tUMPfdl1JsLK20tx0
UaNe3BKK5JPTRuYOZd9ToiL5TRmh2ksetehJ08kdgylVyPZk7L0r1R00E2G6eFBC
ognRpu1T+ehZZ0T0HjkjNcnmCBRDjuJ7aTN072p002cww3FWuVWcSVKrx/O3sHe+
1jjaWRGyO4kUh3F5UJk0hVF4QqSFDgmKUpvnHECduO4fEP6910iYcxgOgcJkJl8X
khFo+sDEbPxWRBeImKpRu+Uw3sdFQGmDz8h7GePJgkkyHlahsCnO4tt7sFnFT67R
Zko/D0JAd5XmtoozU1rFssQQ7uVDI4C4keJ44dndWy1THjCKDFzfxxhJVKg2XCz3
AZ01OH6szL4/Eoh9FVgpEaLL7KiuX5sa1fzkd91AJay4hR7ze0J9BNfwP4N1QIvm
K7uKyYi5NmsIzxuCRMZM9mzxt3npRoTARIuOUSyw76NbonlU/BMNfkN1P/p3xvaT
5gpNAs3mx50HMnWULGpMMAH2GfxgwPpOYwWfcrD7TTwBhGRxgDn6GqJA4u7idMep
2UThajVu7SOFkMNVpoYDQic8KFK5u1ZYiz0ixY/Q+uoqqEly9zttjhP/0Zsqx2hf
oQulF7D8sstB2eboF1jJ3hKGRGV/s3b7P7yDK1QxuCUJfhu2Gpuge4vCL3OCAJKQ
foTajwagzK9Xgh76sc3YqMmE/8hoT7gAM5QGPjHRs7+OlDtnxH+0Xo3SM8xtT7bW
YdRRlC5c3FmD0dc6N1SjJh8+hXmQmGDAVi1ab6qSXXFuQozdViFbQythAJpJNC0j
pQnDlFVAR05uzQ45V5sYhBW1pdB95N25Oy4YM9PB6PqalI3l3pmklfmbrMvHvtjd
EpF+hJHnn2Xkwvnxv3w8qLQRRhyIl5OnBrXpHHSYIPucrlYwcvcYWyl/G69NlJVp
egngXt943OluE+htG1Jp1dhr0or4HvCCvffMwpB0kdaNKmdlbHf6vUpNxd6ize4J
RaUTfVysJ9lk6TSCjenN6QhWj/ab5ille5MUjAgkVotm9gkSFBWSMI4EjeN4NSM5
efdXRAP5wK8nJXGtFd6Jju4JrA6FO0Tr0l4ptaB/Y8lbEAA82sTyuTYsaGaCVGso
5fGMltouq0tbf3HRNDbk7PuGW02JKSWUiKSxhr4DVIObQKJ9O3MvMxz0HW3aPUMv
rZ1fOj5JMakW4B3krgwSsU2Z+m+FNZBuCep5tRRLr11fEHjalmob8MEYC3aWM25W
YhrScPGpFxu6pwogqIEbjHXta2iBd7WcgDl+hKNj4C21DkZLiq0sRAzpSM/LsvP4
pSesvdQ/HwNRijLe5uoYirPz7P2NKM2Xig4Xe4OqNV8TY7L29nfQTO9l4A/nOP0u
DvNt8evoPu4XvMlCvPnLbjCcyy4BVzc5PMV9ol0/W9bxyF5JSXwuXDAXkghbSzQP
LydY2WsL6G6KhiDsng6Ue6+GgC++jRgzLkeYK4k+4b/ct37eemU8f2G7S9fBI3RS
PjIYloWznDAzTKejdZat7vW50PsRaMhMtLJ16CP1R+/7OEgQLPhTNe3k5Kdvmxcw
7FFjiQwqNBUbEsQaX3P6FeAx7T/EPk5dgA7U05irMXseuzY7s1RFdHgFexrM/OLm
/ff6y4afFZswzLzqgKWQjiwuXOq+RuSzULxH459plPpGDZPe50newUX06AKslFbD
vN1MaisjXWSmiVDRqCE16heH3lGwqpkj663gsp5dvIT8E8VLXlGtnNJNeFO6DUMA
zaBfUJaThUBpbNe1lo+Xr9HET9IZiI24eV/R55ISiO1jtPst9eoJc7iU6f61IJhF
hKFapFiOAmhGEak0jCOs56rHS+2qtgj2dDyoq1hSQpYl1ZOtZFtCglwHYN27NhkB
q3gQWBkQUV2wum1MvEYf5zSKkkaA0N0Dx0m0pKaYC+mDDp9wbogbJ9Iqryy1gguV
HLqC0rATzybm0fYwPgQcfB0tPvVpLzToHxZi57ikY3w79USVZ7jdxIfcgrT8jqz+
zagAiAlVc0Ja7D9UnNu8NmYmKThaHZ28CXH3tiCwcD9+50lK9YQy+Ra72wTmMfW8
xrZPFEAPcV6tH+M3tSC4nApDYnnBIWgP81xgxvGA4iHD5C4f0wfIrt9spyrdw22c
eOT38FrXBYqCSd4tEIck5r7xaHBjmK5feBBoG5MI0lucoGf8taTwIgnleK54NIEv
SzZrdc6vYwrgyCUp9OahBArSPa1HLjewuvxcsg+S2bNTC1il2DuW+FVoStQSLEQ1
jHdfuE5BsijYewEt3LC0utE2Ztuj3stsbrGwvJGIbTP8yCmLQortD3BRP5epxJZG
E3fQPN6paS3bh+6t8gPTLXJXPNPVPbogMZMLoAZQDpzCL4vklz2HThharcbRQnM9
G+JsjXgtw9GSnSMnwic85qvkysCGPCD2jQOHyV+Uf7ZQjUhUmIORrnw8JPS6zw0i
m8BWgP0ERoTU6rnD1MijeToIx1AG/I0VhANJ2+MJQlMHUia37Ocp/YHVhgLsL/NL
0jOQpMZPc89iSwap8ew9nu3F1ctOwBAi6KVbv3xmZUVe+akK6Fy0BYK2Aj9+HzcK
w+WzxU/zu6wyN3KN5dpp5toRvryYfJQuqMFygpjufF/SwAdXli/Od7RP4gajxPPR
L5yHGF/ddXI24XweTGQg1zLxHNMoQS7gqST55Qx1qCUJ4VdRU6JbQjSKzMMIY0TC
dh+6gnZOfcZ87fHPpBETI/L2IA8Rz8nwr2cRyL7IhVlKC/g33L7MfA9HRG7G+F/p
TbkrITmMRfy4AJHD7st4OhvVheKkWMlbYo4y9t55BViVB+BaBTuNO1kNFQbCMV2p
4iOf/BlQbvya4WOLesd2dN3Oxluh/GmOf9aRxYSx2FTWFli0xce8i1tgj1/FwQUU
d/PY/zw3RyA9UfvOsuSfu2y8HAEAvViD/UqU3aeYuT79hl75u98fqwiTHvGboaPI
71mi+mt+RqlwqE7zpszM1VpFjjwfABfMucxIYUxeVqpHT2fJwKPMUFFjz9+KvTNJ
YsSJRjetHsWEVEb2J7c6ulEm/98ew2TFt3xUZRG0kGPSWTfdkDAn8JaeWn/T1lHB
TP1VLazQtUxFKY2BOgKOehusEFQ0ebT3xfHS9OkQFBZIQRi+JWvKDn0rbiNzOh9C
RKUQvMNdGjgszwLgodU/Xe5XEfdyXRAt4tAzINMcESGguzoVlbaApxFGYYGC8j1C
P/bUZKb6F38ejtKz38zoEz4cOIIYu5dClCoKqOpiZGLet6QnOQdzyEBHhL78VVfY
lhk76wHNHoWesFp2rXVIMUwMHKj65VeiWxKeu6+OPv1VTxYPTZi0m7ISsbgsIX+Y
FWVL3gFcl9cnSNyFHuD8Zt3c/VVxv6CH1h/IBVmu1dkOzj20XHqmi7aJZEM55A9Z
YrN91KL3emaD8voHn1V2L5/a6H8MlkbOGKutmg6doEWIwRxZgtZuzvu4DNayz5g5
zG04rl8vRv6HDrV3TfvtxKBqmt5YFXDv4WKfUxSPsWm7E/uFOUcjGa9azdgfkNNB
ooDtfty41RBqncCgULb5syD1uBOuArVyGHvanafSJ7PALh93Bjpjr0cr1y4tCepT
sTPVm7if6/6xO1C+YabvPuYRZLAU/6COk2aUwBevO9R1mkfQeOW6+tyXR/mJnKGA
QoN4WJOnnxId3vMt3/lSdFVx9PRgksaDD3EwCPMjUVIxbVNlERZiztzp9YYAy76D
D605uVBkaO/osBT4WhnVLVRrtHQokzGjqQRYu8eqRFX20mzxZLBiCQb50q09E/El
iubhX36+yaEuNpxZjcebuWChq7Dt8HedQqt7WLG8nK0r2LAKX3whzpPRJD5zLdao
bVANOjOA7m3iY3a3DTGsAhyiMjF19hAu55HT74NESWdQbxlLZxD80wwzi1qucuyD
7O81qrR6Z27d1Dt9tB4Hq0qKXH4xcKVFmjmhkHJpLI3AzW2f42VvNcarVSaWicko
SS9jekS4bRh+OypfsmOjCknOY6DCFWY26XZ5g7NdkdzmTNJhkkUMwECT4yNOacgM
fDpjKSv7jX36/SUsG44XCdm0PS4wJRxzAtBrxUr9nTfkuUt0z8MgVi8QmL8Ob9pz
bYCN1isS/xhKaooH6654Ii17oyXJMr530kmGsNgNlDcpTPSzV6ci8Fho7uckVgeQ
79fK/xMDPpEB9RQyC1amZMxtIywI1wdY+CRGVmODsoukpABvNVk4mxyJDlUQAPl2
yWLR84xR4C4BYVpKko35WLhOn1kl6TREgZmrj54D2nnEwawXMhTdLVOMeKHe6HaB
GSTbJ/uQPxT7fVj527XkfX9VYsnbpp+MehxWh11olrd3AE8Rb34vkzShpkA7Jyo/
vEy18Tz9MjyUaQ2ZcxZQGYnBiQXEtp2NQ7dUAbG6s3mw3wLJrvS4Xh8x8DVx00R6
KLH3qcSrtFvSXtQO6BoAWTSsNnJI+sWjQV5ZScJI20qL927Dw5QZz54hA98JcNh3
o5XziawP9TqWGRfaF4MHoUD7ZZr1xdF1DEedMc6sh2t+vfWhiYO+GC4/ElcRaAbI
4C71jwo1XlcNEN/GBsvP8rDfgCFu9eWOyqwniLr2F3xCbkQ6JShRxPt6Nge4HyUi
YA2bxHp2Ar//8xq7PhXMI9lCNCcYXa5zOrLM+7qgqWqLPgKM4jwwObFV/z3arAFL
I9M5e+orNKubHsX+C2bmUWPi76nMqYQZM/cTyJ5DmLJGkBB8OlT4ISZ+eFqgrL+X
1oldsf/+VZ1/Yrr1QT/CSk0PxyydhFk3d9ZAh8WEkMSytdLnRICpqChx4PYgLziZ
ZKg2CsMyy91YlXb3+4sWb2+vqd7gqJ/AjNmI/5YxlOHxgpeco4P1zYlX21k42so1
GcX6VWn3zIGvSJDlK+R6iYrJ0N8ut5aDFLENtLidti46rBmiOkvLFcpsK2HQlCEP
hYileGYID+EcvDOpl2C2ntfyVjOsYOQBe6ySkKtiLE5ktf3cst6HYj/dcDHjwmkb
JtEGRchEA+zkfWH2PCJmM2/IeDGM6mSj6HPgd21TL11HRkAJQzubAbQzcMiqwRfU
D3MyAYEszTDmVYqWb9IiwnR6MQ146fKk1qXd5UDjO1okH5Rb3dRwNt3yWjhaOOhR
8Ti1l/0o6xkjn9SHsFtehvEc2YjaQ28CVocuCMoRNU+gxLAPyfqm/X4uDzvLnURS
SU2XBNJ3O/N+2L79ewW55zR4BzByAv70fvjNhaGoiW7iLG000gOVcmkeULUtXWJ9
bDxaUdae9AkzMTISvi84oEzD6CNcj4SCC/RSUU1QiZsUHj2mx6XOTPMY+dP0gRtu
vi8NslsR51t0iihCQG0dH/AWu+Oym1tgfhVfnkX5BAyPpQM0vLh+fHgkbfIiYluG
F0Fr5JDx/RE8KACG3lcarnY80JfYIxbXkS8gAERkZgY4SAl+Uh4FKrzPF/Mu2l0D
H6pfhNnrhJFV3r6oIXQwvIZSxm/jyWeLQ9X5m66snY1FlQd7ViGPRWFyl8swbysi
t5ll+FOs7w2RZqNxAJ+GrcTivUlxC1WooByPfrHu2nYP6DskOb2kgZCf1jIUkLBN
BfnmyAl04em5f1CsQ9pGnpyz6r6cGGbR36xyZlyM8V7XIvH9MxQPtVCUcbKI+7+a
7ckcRqYXdZ9IT7Lmi0fhzi9lEljfi7azkFgdV5bGY9KorePbRL972xISnAWEJ1YK
3W1i4UKlrEox9/y7c88PVLhH5i6OVeZAR8qBucxRyNiIQfp/XQsPpiT9LwbFNQee
pHbsags+PQ9ctTT6i6GRx6BZ1BMhkJbNkkAcX7AL4SGCz+QUVT+twFe3y/rQuoiA
n7e6EvGJTPo+z1Lve5SYnCsgQiSTqcjPFesDsfKK/zCJxZtrbgmLASN6Ex+eh3TU
CSjNbU178HWlruw4x8WhiuVAFQHZ1gUdwxLWYdp7g/IwN2AHIuNbNtlW9kACHFTj
ygiqZjgkEQMivDjYBozeyZdExRx8DLhOOM9a24NMiOIup/O7XDRAHjaiNTLjYLP1
JAJzFRDISS6MmwBoMch91U2ev/L/S6b1EEQX4kWXzFltCzzbaxq4F4JyHqt+FUAc
KSU4V6LnK5UX4T4V/QsSPCSGnMcguqWbLeUObqIuSNY4U7O0sAFa2oF19piNM2qZ
J6GhB2CmzxTFd1rqlCz8u3/suJPbP7sFbvr5Un2V5AQT2A1azveeKf5WGhb4ST4+
+8u8q3drHb7Cb3zo29P67GJaPbOxxakh83jIQynEHUMpX1c7BA5FkeMW4SsT5mW4
sc333khylvnPOjrajSDJpJv0pYrZE4Is8I5Hk2vklD90V5CWI0CKwFRYOTJoOmct
SKQWWxCjUAQmbDu58eaU6NXHKBx3B6CXTh5/VZoLKwoTnSIwHnKStQihxvlRMaId
0Wv8ajY9YxXHV9qnu6YKU7SmgHfLgX8fEFzv4+zNcYthuYsyBj+Trxq9c3p64D2y
pp5Y5+yL2xqmdXBAUsqaElTKj7stiApatQDGzzDz7rqBOg9PNwIkAryW2s0egFLp
MnWVBDK2Js3TdEejWjeJKzsW2lKG18Lof5EH9Wlf1JBJ0NNPTUKFi+CgtkhAcDd7
sMvP+9nnNWU42iYVRIFGhqtIKWB1+lrZZiRj2zy+XJDyD6m41NZi9jgnPIZTcrCo
DH+4w7OCprCjDtL3667+CTUQoNob8AXkrc5aPsA4B9679/kcwOO9liPjA4gUA7JB
RuDBm6TzzdmEUucyOTIexvXjFmO/EqgQcK0gz+qYYXFD1zm1CA9LIsM1TlCtw7zx
v/VSlhyhrwG8uCg0ALXYBCJ9RoG1tZzzPvXVufHS39PK7FZPIyzW25LPLfH0na3o
vpet2C35uG5q/OogLfiU8oIOOByrn9lt7erPwU7oZm49K6pAY3kdyRNA1LZiDAKB
F/cvCoRVbXRXzGHUSceV4nX385sJApLx6oMfMRdZPTdZXAVrFH6v+8IejUYVnKPG
RjX86SgA/sSa3Z6Oa0N6c/w1KJu5KiN8EcAu17dqVb9llficA3uH2qefcX6Ufx3N
ZL/i/mu3ggE9QXCYdR8LjwEQ68OkyC8U3tunP/axruZvIOXIcvIE62yZd74fvMlO
zUHCnWy3X2woohPZpx25Pl4LfTMAyNjGc3yeUXDGvTgtpZPnxHeVH7HqH+19rR0m
sj3yGPv6GJWfPz7+I0TRV9hnEz6ivcCzvarr6p9oUFkn7FxuIRj5ImUWn5txOobw
JziVJye6PnSnJz+7zRvDp//YETCTCBNyI7UXCwwYBXhKVf2WjUE8zzFSZTdPUg4r
fP4Kwkc7WoCmHwCufVKC2H15K+l7JVH1c8cdREmqELPXg7ONiVjVDZ5wzbNlZjY3
0eL5JnSdFXcmVXncAYsTl8G/7+TPNsVeAHh88yhsaoaWbcFKKRVe1eLYb2qkIt/N
UOV8dzChqpWDuVnTpN6AXgCKnvZ+Sx947W9nl/KOIyhLez3Xdp3bHuyeOmPY4UjC
UtSO8GBke8FAJLX+sFMqUDIUe7OEwBz2JJVhn9CXxUkRFXfMfDG2ZhkNCmkzimd+
eaD/47i7JV9nTzPypOLVUkrHAKTI08HESU6q+JZoDdUM1/VIc5TlbCefcoBPP6ec
W1fAzMDKqaxmw1v2iCbfKM9ukJWhLGVSaNx+A6wuMLd6nkaZz+LAHDvK8Biy/0ad
0QM2oZfi0m6qtMysMb5/NVBwOCi2qk0pxovbi+lTxHxPD/wJnRi/GkroWEEHAxjN
e4vRZRS/n4AWdkzqpImv6KHGOOQi5DA9X7NiyrxYtQPNO+eJy9H6jq3V6omhNiU8
z/OGCZS/f5umEd7z2aye1nFY0gFhUlHnPuEKYAmTdZo5LhX5LaRw/Hx656ecV3Wx
6VQQExXARtkABw6Ya5aTTTWA1O7f5k7XR9XypBoA6RPBudjPGSf3AG9CeS43lR+J
IVnKXVztzuurP86MFUPJbZToibrp9Z5YFpk8AYLCJ1NXCuECQvMpmpwIW641ud0e
5ISHqrIObKsNqXOW7/BVdO1bRK/W+RZ5NL/PPl4C123BC5P3pCPGriIPsgkhd2Xq
nJzWzXwiYT1jhCQtA/iSNXR6yrU9o2ZMW625ri74q0HddveJRivyif6MJe7pIBF+
4Wnrip+m4UbEg4PTeCvV7S6kS67gTxSs99hssHsNwvklPPRWWoCLHWdALuvHJq7f
ijFV4y1ramQX2Ksx0PxUOaTUJuD4D2/vQdg68aq9BBX4tbU26m1jSzbJUGPAU1Qh
2wzxKGEdvpaZ0fjpS0T+1BQAOcN8wrUp4c+JEuCE0ej9cEuC+fJ1fY5Zy3yMxC54
n/k87XMaIuF3Lo8eK6+poEJYfwkdKoZ/LM9Gu8J50kSou49iuqGxstIcEtORGpX5
aERKSziRcFIEg2cWf/B+ErG7NnO3k6wq2cx0gc8KGZdcxF8DBcPekVCNVb4byspu
JZK6j1wzK0Rn5bqxhta1rSWcXZjTcTQ0pjJjdWcrpH0kOUx0rRWrn/RT31HbUHdb
hUrDx25h1DJ63u7N5iaCAhglt5qXac95H8s/fUF8/aEzdwyn+pE/xE4bEUDtgUfx
xzNezIcHlb5EAvJ0YyS6S4ORTI8JOplKKh18F9gz6pRKCG3rMnqX4iVyd54sSOLJ
GGOpPm4asGMeYSXg386qKbdppHVDSUbiHND4U7ztdLIr8dZfl7rRk7KryxYm6F9h
FgWxt1DDwVGKeYkxMgmToqGPwy8hjtr7cXwEIhRxuXpVMqUnWb7OpWf8r/Cjikfa
RZOYJ7BJMbtoPXLM0fwqqlP2z6svckcM7PErs1oilqVmlIKCFYLe5m/cK1THQo3J
5JpftjMNXAtRWYEIaaJbskZUyNRGjQixxSleDX2sXf1qrir3fLBC+atq61gYl0Mj
WpzOMMw2P3dRWJkQyGY0pfSfqMRR+c7WYrVEqm+BvlqNehKWyrq+HS2WhD9WxWoM
hkrEWOYsP+ErfMWAlTFx0MdnUTdkFjdRbOPDWBAZ0yOiLCIIoJK1vv3sTcMil3Vb
AQR85zeFyHZ4GlNwpX92SyS2s38B/WS29q20VuhLOIAfMjZR1DuaqfLUkczRIJ0A
k6h98yCUB71Tz1H9RedwwX5bah+RZey14sYCkalTG5MujW4V01zU08TtExs7M+d/
2TvQvVcqJ3MN1pig5aqQ8KMaIlk7YyhRzrW03YVDZM1QU54dGqh8X+z8vTzcei7s
G54lxFSQs4ZDszp6sv593iuTQWszlfXHxAGOyc1YBkdkafDHUxMep9/CuPCaMSss
KaLileoUmMpi3Ig9/M8mG3zu2S8Eh15d6Np8K+UohnBxKGAXwXWPrkuKoduN3fXH
/i62c0bJZ4xIygatMwDI6Ufgj9SH9mFQMtjTuSTzew+nr6SOswVgUAT42OSMy94X
Qv0T5HvU+enebXAhhOvc0EMqDKGDhRu0v4Y/mEAEdBrP6PioTlzZjVUh/EMSmYFg
I/CHzxJ68U5LoxH6Q25PApRmPNnxmDIQwmuF/4+8dqjkvZjfY9uZ2reoAQONOuLF
vLPuSO3MUlUVQEJzpd+qGdLEfmLx2apqHce2NsfwqSGXZ17ZDb0k9Stoer3nbf/g
aFGbvuSxRDS7XTmKuigDJo0xxTG1E/YD8h0AdH5b827q2Uxk5PbslRJldyaKV8dj
hnejXSyDuhsWcntln8CsRqbQg3Q31oh6qOoiTFBZxRG3nZSaER83nvX/pRm9klLr
C49IOqtxDuD86zGUaCNPYfMav2AFf/Q53rt9xzpOLrIX/e8BUevQExmk85RHWj9P
Voqt99pKBwDA0110ZRONSTC8AMcZX2wp308pBQwUVTAr/fUNy6T1rWwuOwdbWRCt
L5vFCfEIyy3TIuvIsoQTLhnZLvM1h0NFsJsrAPVEfIYvSbn6ZHn115rN9EZrB6x6
prU2nnSOcrh0AS+XoEvu8f4C+gMAJIpZ8WGc7EqDFE0HlzzHFslcxemgOhSeMvUM
2EHx8Wcaio69UCHdMMl8GprMyO/8c22uOO1DpAeK2PYci3hH2mG7MxOHW48rahol
WqfhcFzLmMjkJegj+yYBmynv/mb/P8efohTQwsU8nZFYutrt/3aRoy0nrBe6owM7
p/5QaYzU8mJiv//ZWCXlbBKRRULviw7/Qkci+8wOFIym80uYv2ae2l+0iBfMTzCP
TtCYPb5xTeniAz5KNBPxYoXlusxtqSgnLB/QkyAdXxbZTsrLoDyXOIyNaeEbkkPN
0cd7pIE1HBXjv7nPWpb46FiKWhjibRvUjdwHcFqOYdzVlXwmmwxVlJ29KD7elKm/
+5nRg79pz079Er4CPNk2IltalT+YOil2cfoUlUST3UcHP1htDENa6ej+uiseW+7p
/g6TQZIu/ugAqJ+p8tW+kB4d/EG1TMyXUXs9DR21G0rC+YQYPnvQfi/1920SDQSk
HthlvieNiBAYwR89Xr0N4BmtjbAK4kpXSszqaoiGIj9WXRDATtvY4iGA6FgFuC5E
SiyCXztVoyeZzMSqufJRnxNPup35DTn4B6OSHZldoFEUlusGimdL5cOlRSk+W8tm
kE32WtLtdttHMX9ZpgfrRbnuOWHoobSROUfifj8iEYcxe6A9Xwx3ztE4rnmX802S
gD1sTixZbF/aqFWMakK086CBxjqQDinMm+efjzqTX4x/2p319goB+azKVZVP9DHZ
h9HzT/Y2bSm/Gl0Ubv61v5rpiYUXhKe4UMc8a+wehv1LgZA8qTwqgCyldZW9xA3S
SKMJc8X8+fKxFWWSjJqaF6wm+aDGVkCK7M1B1TUhq8u4MTVNJ5ysJ66K4r/eKy/e
7Xt2q4+eP+mB+t2rRDp9/mqqw67I6fiDEgjNFcUl0KRiuJlyIvTC2G3OX6cyOBeS
9vsAk12PbUnRdvm524WzJznv9UyYFpLmfLCkkOFjHy2ISbvECjPmrhgxQZ0zY0In
kHyZ3AhVbjqhQlBo5lHyWq3t+O9t9DLfHeR6706q0Q/39Ks+d+ITmzMzzmw1wuvZ
pFSesT1syW22XZq5b4gBiHuQFOjRbzfc7al5kTAxkkOFhwuVtnz61O+wBdUy5O7R
oi/zTQs0f1+LgiMOhZhoMBxQf57jghdc9jD1bfJLglblz0VqRaVX7h0rtszFdAAE
NF0CXyxJt16bXhSGjhqoJHTkww6QLHAalOsrgi8nj9nWmGpG7rpHBMhNpkXuc5/4
Rus2yHkgEDFMWlDwIIQK3SFhqvkaTocY0/HCexyndHs99rPkpcqzoE10qXzKjaNB
T3mCYR3DL8K4pxDrHkV5dyalu9opEVGK7KY/CI2X938KMWwRmwyvjohqFFXBuIAv
W5n5MAQ/r+Q5igaOr0C0vKAmIH0WAtutySGbdOsWmbT3Xm87zPfUGU8+ahbCVzsO
M7ZkSTIzLCDvY8Cx8dqlujZeRgrxvyJ7NFhzVliRuolGjypbIfQOROhAbaPnrvYJ
zIk0JQTOMOsb7g50HN9vaM5p2sdEnTyy2LisdkR0Qfg5tTh7b0tGu0GsNqA98R8u
H9qW/jfm4ivobkg1+6gm4b/seZUZICm8F7UBFqTOFWOIzzAxALiTsA25KttOtAzy
SiYolzAyKMuc8/zyIQC3q/16emGN2XKYVH7JLtUzf9sqErk/IGOdXKWC/uyrPHS8
5WevDlJoOSFft/OcFFEmuWecIr5voUJn0J8nfqZMcLf+0RwLaqKwui0/ZRMPou7C
K+lZHmaUiMv53bQLTRsC1BPbWpdYvgwT3A19xJoC6UPRrapyN40zBWuWlCExxwpY
w0hwzVAMlWcR4BdXzboa1GoAouX/eqd64dw9EroAMr6AJz7a7bYFMMuacSKvn2N4
VmSHwNlBY7zBnktoZEYqtGIWfDCQDJxU/D/DijINDhIxeIK3FbfC7OjSprPl+A5t
lzZ2pbvbEx2ClBj6Rr2yeROSiSo03K+RuPLZqwMD5ACWohSQgQHnWgkfGvi/GyC0
Rhm6rpaMZ8KF47kSu9E4/3vG9LQ4nEX+DqZTS85hJZVGiYDELKxRF+Pal7K7QCQg
kFZvGm2S2Lfb+Dsn0g/ko7iHDKWHtC8Uvw8l2GhZC2E7D8YuKt72YOaVSG9Ugs7g
lrh5Yp7ZGPMA0XEkn26WFoTPiyQ+dWoWkOT0VIzHMAJXxzU+pNhDf62j8Baf8ph1
rwc0uJaShmlwQ8n87EqCBDv6HxNatGY/1nR715gxT5uyfW2nDvZF83XfnOLagp4o
BwNXGrtOa3VSRGwm9JqOBN1oFACW3OVnpMxw7UYy1y/6kAVflsZ0j/bYS/rVuwLv
4vo+DNXZxksvoi6alT5ou9HEInKxO7xDlUS6yFdyZOtKENtQp4z2RnxoCjmEfSmZ
VFaYpyzXTLj5xD4JK078O/QVVuEFNxonWxitgPKJFxU5m/6B0PNjBQX/LhYI5gSO
hwOnpKT/PGJD1aMFEKR/cwLQuYKhXvyhkBZX5C6iI1bF5jVzefrpdzcRLnCNSZ7w
dt3W1jGOKEt/K4qsz4RVn4+omPWKxKN/aQavNPztzShtKa85qnMGEdjJ68GoJbdM
rK+YXJ+pMCpFGm/G1Q14lbAcg3OTRnBPhpBit7dTK3JxFr1zfNJIb+tOCIhcDuSV
IeE/4d4Y0k24ymVOTUSzPhMB7tx/IHoFXc1f9U6uTUxQ758IiP66OqucwB+1tOY3
XUISlMuwHYtoP49uvzxuDTtqklEzoxcoqaSKGmwXHJcrAj0jgXtkXWwSnUOYY4vN
lXR+Aqvl4Pe1Qc5lmSc6qHJaMCfnAEtlWA6B6IvfHFQquN2HLqym+Vo3o39HW5N2
hdpgCulhwqNgOVw9i/IVExndX8W+VAumZcW4ZDNZ53enWapqpGzEOj7dUlRCOKlq
IXgH7YITrM0tYlpjz/goAnL6HeAkF+C/XS+2OR6EKXCkO7fiWcGZXnjWWXmH9bhT
H9z5ATp5CE9NrK7+wyOCSQBvs0zDfmspPSEJ+cSj72+YsnOpZRalWI8V0ZSfWmfW
Nxz4FW6YPDs6Hssl6l3S9UFfZ9Bh/OI5+RXYziOpCc8PG+SNd48qkqXwTQzjpMPu
BTEo6SVvpKhe3qdzGePFKOxKb8I7dxkw/9csHA1HkcM9FuCFZvF+gtxIdc9MNL6g
kQF85kZg48oWVnF1LkoYZ4DsyP8SMARamMNGRIIkV48dXHk3aEwad0q3OvCbYtpQ
JIOqVJki2zq6tF/svhzTMyAbtkpcwxPzWdmjArlamawn5Bj/+z2K8td1IqogeMuR
qnZaelV74pPjY8Kv/UWKr6h37MaUwj9eMQe8nsgzba3axiaPXRRpXtll/b0+P37g
uWPsmMOn0dHOZTBnegqxULYPkXzKcRXnMjdTvuGdvjjJz4wqrxLra+JsBBiHbAMw
RSsxSNzcTd/HhvJQ5MyzmS+71Fvam5YAU08iRWqMEu7UQ+bosJ9Sxdy2EM1HSaUI
7fd/GuhkYQU7lDzUXPcG77qGFgVINZPfHtykPJiW60dl5KFr8R5hd2Bo6nfDQcSV
bJamvuqQ6i7Ao65seOwXYUFRtOqPpFHKj0sCU/B2f6ZDnUWbeSDw8LH3qUTFqX8S
ohqC+0A2LSI9WfTRgMIwCHay6HepmcYKcIhBSZ00zLFxAPQmJnCgy4Khe4h1ALzM
Kjj9ZDdHIWvX4UzzgMw8Mz7U2KhcXM540zsVaJXvbhP+CYjy5tS6nOVgmxi/PSm/
mfIu1LxfskEVexiNb9TjO/JQYXUzmIbZs+MyYZp7YJ2BM7SdX0qGyU8JhQZkCgy9
KR2k6AvkUwQYx0weqf7K2tFw71j57TWn9sFQN9d5z1sfyY4BtH2c9rRNkQ/zprfm
w2M2GOwFOlfjfa0C/sJeatM9TM+RMzAoXcizUjOZkITZmN14lDcP8mOP8o5+cufz
deY621ZiyyTRqo8pMW6fc72qFOj6P5sayY9q5Gw0i/282sFVYddYrc64hgLqwgFO
2x7FGZelUTskI9/VgtnDNQIg/Mc47N9ahO7esXB+/f+h56TSiz1FnrSK9Y7lOxid
5aoQ5U5IHwtsRKZ5xm2T0umHekDplCXasGCSyjvdi5t8JTfzlpHm6OcBqmyVnCFo
vk+F5CXc/DHps1f0nuRbSUF47AlShc5+x0ZjUUejrkg4TSbjvMYnXyZ+OQuZXKrC
Q/tXUzLDJRBA9Ew+SdpO4GFkcJtsE3nC+EYunGWTSCYD3K3hK71Tn2525oD403Qo
51utMz2dGLLNqFfj+oL4Y5UY/1D+fpFqBM4IJz8Ymji4AjhBueBD7QaSR1TQ7RuD
gZLWQXh3YngRJx1el2G2nj8zm1uGBlQmPVI6k0uQngIiXV4zE1fGmiw/1i78zTJL
G94RE+0QgxcS2tUc7ujLq5dxNpy1+XTE5jEYBkmx0MRSDuvNaqpSNBdzTVzEsui0
s+8qfha94izubi4qdaE+Oc+oc2+gDmPHhRoj7wfZ70GQ/Ai5c7tkkIcW33C0t16s
z/mEYh9TDjDpELbca0GkZFjV8+HeEPTRXcI/woySkcfkRBYB7R6hdDo/D/JueX4w
BUeetHr4Z5NK4O88dF7Dk7mZriA9hJxEzAwR3hAjkee7fTCjtS47ekeQrvsoJnvc
I+2+SeMgFQYlRu3FYDlTGKPjuQ7MDj+yDWrVuj6ly/JugVLZv05F5BIt75BfolT4
6cexg/YlzVYFa7qhFAYG/y1JXmeJ8+yjhHLsd0bN2/9eliNu8A8Cc20KuNEJqtus
I1nKK2xl/YGIXcPaZC/KuxDFn370iNoOBk2IgMq5hPkUjVxpjt96Dppi36q8uu36
iOWXU7iCcGz13RVssz6Us9Ly9HnCn67jCCKaciEX1uk+psY4V0ivKon4FSC6rZWZ
Q9fSmU/+Lqfa72oG8PsHAOUCmPWU2saC++VMGATgBbmDHutmG6Vhckw+JViIryeB
3RsWQ1gc+fOZvk+YaQZd5LdceHF2KeOL1QiF2mFX1kHaMXH+2L682pdVQdoK8jB/
vyuvrPxRCdN/+hpxc/Zqm3WWXj5BYDEcgzp2nvGr34uxiDwIPOpdCVGZEC82w25G
SAc6z6dO1p7rmf+sY0pa7Wq190VcZxLR3Hz14GTlVOzK15nZ4o/oDKUhmMRjm9E7
t10OlyHemSWGcDsBLKqi7wNH4wh9tYQs4oILlItRZ20wv9vi6bIQExYCYMyn91mJ
dP394uH6EoaWXs0hW1o6i/82bAw2ZmduajzGJhI8FORYBSoTI7E+7T4SzjXJ9BCG
8PhXiwlGQB9gJn7CETPfUkJh9i46/Km069MrxEJ7erqzcnWCwh3iSzQAhwq/GmZT
aPanYg2tVP5cMIiFKgg3mg5iH88mTnMEGnv5a0FKmGMWIERO4FuxV785+aqZBw6Y
xZvdftjRwefOlikbaYFJ1nZDeswesQoPZ1W9Q5640JAt5a1UrF2aP6ETCvxG1eqd
FE+PkBGiBH6RFmk8V4hrhjnj+6WE6CupXP3Ox/39LUIHeld2G/drOXORuaAU1V/f
T6NKINA3aiEjPDj3t93rLgfK64vLg91PrZpsC07RRM+KiDmcos1QMTtwY7mkuGy2
ctQ6/xdg+BaSyGUlTHdzsFpTrnBIa+JWU7PafJWbtyQWZP9tWMDJe+zD0Nnef6hQ
QEkQl3F99VuRgkfApcW+y9FYt55gylFdD+FqqGnKrtkBjCUU02alnMxzVX5nJ/8d
xkgc5gAqc4kK/f0DkqqE1E1HT3xh/HGcLviQzdJ+b0qkoKHqV4/zsaMMDY0/0Z1o
dGrTVvjb8H5ixTQaU2Mp/jRcxZEtEDS/P3AeBWDUeV+b4TPBXLeLprNNKkZ7CJ7x
abcq8v0OCFata6bEOFpMw6+w533Xbm2xe3ZBCQwqiuJ+BLxjSkkfqo3eVb7Kyl1S
2VkRx4a0EYCouyKM6mZxIfWlkD8i6eSylK5zpnexiuIEWAXIimAE88Flmfkpc4Wr
o+c/WrMcD9cznp6DtbV1l0luhPYVVDxtxXgc1VXcMnsEVmor9QT+t2LYp4caiN+D
NI9pWMgCXZ91C5nHKw2lQ+mT/LEoCnOZR1wkGRLW//xNRccJmoa+12NCNhLdWFdZ
cNaLj580veoBg/HCZh3Y7QjtcQnnfN5a97TTAbaYZM3CWZEwB/g0UXMZBqk76/Q6
zvPVzON3P2Th1bzu0narqQ+n9X5XC1KleNjPG4GNh6jUPfhm5ZfRDNjoBhV17OZV
COfj7MdLf72geaK/oKv4IwxYno8FN2GE3q7J8rbig3Zkm4S0pFfjJevCno/WoFWL
bcfLJd9sAe4z+v7dPK88r6HvcYbYWdUOHkskjFoABE9FXtGwpq+BnzAzFcOvvjp0
FMD7zwFs82SZvVO2kSw4ay+x4OEQCbQpSz0VM+0RKOfLj5+Uc83SmHRPDq4HBlnT
hP+3tFdZJw/qtJu8Ns9QG4JoQcdvuj+vD8TGrJ71y9aljwkPZNC1msiLwGoIY03R
8WqTD8VlsU6gKGqwKyO0CuSqDhWP75cOstjzYQ4viQ17o6ir1EIOEyCvCFUqxmbR
Wsz5NMElHY9zQTYQwjfn7dDvBXfbRcVDlps/qq7TSag/TbCXPpJZJHjWngaOpXYd
xKgR71wN/EnaDC4XPe8i/C1a5r/265oInleViqxhjNTplok6ALbsQ2Wy0VvrlfAH
SZwM87GLZlwRwEsEgw6cI6FP1vmjXlvf34b71+mEh0iffHlzEd0LVWQxcZTS2Rv9
RaVijziXn9FrOd2Td3uEVt6/pwzZKOyndR/mimTRmh6pBH46PdTRCjCTFltZIq5d
mKyrcWnpDW0h3R3kflqCOZD7dOI4xQTk/Rz+r1Y+2xtjvxA4I4jzoJ2wRTnVn57P
d9g01q/Zn+isnOwJ+0DABaQylnxt+IvVtKBVWwHf77RXkiEGPksE2d0TKGpEmNFu
Pqeheh72fVhRACgvowdMe3TXTJTic+i6T6/xhJ8osya9oGmFUZgfUYp8kSEuzS5t
b2+H6zIpGAWDfNai+M6WV3OoJLcGNVe5XVjFLawy2cABojTjNAVknRpqpn2xDvib
0ZuN1pIuiNfioUsNKwcwX9meKguXaMI/Xe2tXt/HrxkT3u/5DzU6kYSxEexNJFih
BeXOti2B3VImzIYoBmZrjkmaR0DU88MfbNs8a4tOB85SkaapvVeqRdnVszQgaJqc
CDaVWgSNJsJp0f/j/qBXx0hZuSvflIQw9NCgV03rdbWZRPx7jbgVVSRLh9NpBJKp
cyYgIjIfRgm8Tzcnh4D8I8f+2Fr5P67/5XCfsBLtHGNa3UHW5CBwtrBrfXqEW3C0
ZtEvJBgYkIwD4Z9zzUVYVciAMt0HvB3QH3EVepVz5NEEocwmQh2juJuzH23C7Q+V
P5iX2lDQbM5duobyLwdRNtp8cwa9hGd50zxz5w97ZpBg9gLb/CsqWEJihdXuFwbn
RYGSXWow45kuBP2ocWFKWBY2Xn7R0ugCQi9eqvbJCAG5cJexU4WMXD/XkFD2Y8m9
qsPvl+3sCMTRQhypPUxEXv5Q9kaVYRfZ/4mY2kVAWSCaPFjvgBheFa2tE0Po3NVf
fTvxhYe9r1a3O6wCmY4VqMJ1ev9l0YWqLJzQhZri5iR22/GzrPd81JAP5WvniBzy
IP4TS/MMd9rZfe+ANjj9aq8YoOpAXddZKrWs7fUW867UF0WlmYfy+EyzG9x/esro
+r+mkO9hfbiN9/WoyhzRjNhenrVVXn+T3mhPEpmKhC+uCR8YaFOTUqTVloqVCZjL
7H56+fokQCM8M62I/m75aVBJvGWaC0+wEEnUkr1jedSdOf0iP3D1t8vgqRV+71Hm
XIWvBsGRVXj3T2aRDutkehO+bR22Ww9y9MVzB2yxEv1e8pL74IIhRl/pwx+N6y81
PfwBq3zUDhvUqlz8e40t3DgvKkqyLO4LdWJ+/lBmUarhmgBE1dWaborxPRLNa+Kf
+CADUBjN//whva2qY1Rb4dVzaqMpaVAIl5F+lc1W9N+mo6w682QR8sySYN8OF56r
1ID4MB/ms8qmeYZYk3dIvQntFlvhwSguaIknSMRNMjaknwVGh/cWKYZwdY7F4tAS
4rKVItBdhtoMck+IMdoQibMlV6vwLngqygN4ub97sewJPyU8VG+owpQr7dJZujwW
me79eReGy15y73eOSwLEqwPdQOb08Ng2DYZHomhPYr4GR8p+nfodT3mxnFFUl2K0
hin5o3lQ9vQ/h/Fi1eDnWvJV1D9z5blQGKUxsF22huWSL0vyb1hmTyBAtQLUifdO
vd4vmRmUdX3RNIItRLw7kNNrOUItRKkaplb+k/m14pgHRYEuukwuRl7kTTE1fcrx
ILP03etWiDtsQ+8fpCTA1cqiHTl30fLdW11tXHsCDpntK7qPjMHP2/yNEdTWbPdx
5ZbRlj3wKTU6mjQsnnGxrbF4TWmr/qlI+fvjHqZL9bSeIZZvBvvys8ff6/oG8X93
nJRdgtcMfaw9tu8v/CUnbJkKmFkCt0cc0cAlDduDv4V5456bcja4gfBls/TjoR8e
hnvgHrlnYoMuta78XvgACMhSjp2EtyTQAK/ERkUf/OQkKUWgBfPNtO/jwIOQWj3j
Vjw6NAgQfrg3shuSk87zjBXeL6hCQibx6rqKvHBWYXYNcunzg9WnHTWx8MmYo0Eg
xjo0JeDnN4iN32pyLv+2zcfCkoomrWYkV3TEnLpu0N6j7EXxEtVLRT6qDcHoyxK8
OHTrp5KH4z3G7Ad9Qx698s/ut7uYutWg1jfV3xjfJYDO3dQ2iqPCyXpyqKMnjhwy
n+Qa+ZbdLVKg1G6GmhpxHEkrIMkQwkUlBMo0tlT5Bn0kg48/J7OB1PlUZr4Z/mWU
S4/2RcEb7xTPppBVoKigXfhD1mjJLMBuVjIi0n9gRiR948mwRUT+Pt+gHLdQmsv8
ogkvMvDyQj4qzfZLQ/TIiBM7ROEXby4BOZ3uBLEaAHOB8Ae1sFewr/bOdJNpBfBW
TvdkzlWwGxcJEZY5MSaoAfY1jJXjbEGVFEustC8sgWovxA0bappsUaWQCyz1wrLS
xH7GiNzgm1e9MDftPFFqQmp7BMXPMlqv3pkg8VqtzE5z2j3yt5kCVHPHjKiYEFKf
xh7G2n1DPaqA8JCpMqTdjaGZrQL/V2mN/sfF0y9RuPJSe2l7lwv0696qcfdU1KVZ
LAQChVcboD5Vdut6PvknrkcMcayN6StBDT3ylomO00ANWgRybSC4AQs7Do6RMnPC
A6m7rJAd5pO44MsR8GHhl7J7GjUjg3/Svk12VKiAdy9sosovaA2WfRWNiTy/ONs8
Uh7PSBQR2R8LgajMf6aGkYt3FeqLpXGMI0RkwhvKAwIQZ79XANWdmh5/0Ib2P0Xh
+Fz+0vo88wSpxH0wg4WA0F/11PvjxVGLjgJ3lNW3YlvwXKrh+8kgMmLbjthkR4Ti
OG2UEEQhheKF4dHANXaZcsxjXXZnAMQg+gqzUY+rkm1jEQ2tV8rOB2LYlwQrp5ol
1FGrbUw0iyHD1qwwwXv5I8LqkAQtznl/E0/khQZ8XlxAveqQgwSZobswhtWlFMhm
X05S8Q/3/OOTxVvf34mEqeo4oQpubKDoHfYoxCID0mPF2mK6vlRVW0ydFO1YNXgu
2BAZPQEbFRsUZ6QXH7wzDJZWZt/0BL0229ziWcYWm4ewPG1tSZvjpOySId+t/Y4Z
lWYVdrIqdYwq/o9WcZ7L3gQJroIwUx8V2kD9k9/SI2KsBLTw3wjv9rpvAI8tnMZ6
s4dnY+Hj9+iTPHDJ7XQklQcCuAfT5na8xdW9CusKC5SYEixmsZzsQXhQRo4Oj5v1
KXSREB1PTmaJI2O9siDblFUUjNiMcX9/y9EOKoGR1obmaxnZnX7JRZN1F7s+ILrz
4QPQw7bICzjT1tk72Xgg0zuo+BLYU2bDgRHEvwQL5fswaScyQccoZHDnqMEoMaM7
fIHfDcCI+LrPhXdsaFrxjdTTiWmmAqShrVbWlMCkwcwicFBxc/46zYWEuqenFRhx
FW7LSfxGYtG6MJE/KZCWBykUmQfYjbRY0aUK7+wIdVswmBuaXtlJJu+Dtu5PSGop
2gS6A81uHkjKgPzMUxayEAeWjF/ZNlQ7WaYWrc1v2d371ZEwzL01g5xdhyHaWlUU
omMUttyFrE1zVXnEKc0ENQ+jzTpoA8+HmcDQVVbzhgAbaAu6GhJjTTYMKZw6c4Lw
1GB5xAko/IdPfgOPjKcPjDv3rrLLyvdGyFgJSR4uczyNN9IzeNDANRJuA2Sraz8f
UuoeZpy0i1u/xktP2sIx6OTgjZetqcFDq7wasetUzf6XGx4n9NPWKGuv7Hsm26mm
gUURQmlEIpf+aPGnpbHjUZhXJk8eFfR7xTyfpyOqX7dEKOhSnVHMvanJC+4pz8NG
S3e9B+6XXgftB6mrNaMUlzea3+Yq541l83qTsgNv5/r9P5k3Yk64ey7hpml+S1SJ
/OspMHvqvyD1EpTqtQyzgVqOWVUqc0gBB7+563P52KLt1fyojtY19roh2iJjJQk6
gQJglpGnm6GuQEGOYQ8F9xR4Zu0uZcDrdXnjm8onD1HPKQslyABCZwIf7c2qgmEh
uNW4TyufHjOo+4VG9ebQ14gzVJp1vXuR1WEOP+0knfccO+7YCy5rvL7yRdnQE9lV
Fbxn5Q3Z66cY9QqkAfjx23BaBQ+lWRVCe5risInimd9gVA5uTV2g0bxHxx+AR5iN
39VVyQ0uYhw5hrnwfunXyrFVR+kVjtqu4w/rYbtuYwdvsNu6hi2TOe1DDZ3rADZt
dPes2TAlKCyHStSP3kE2ok/mYottI6KT8gC/+J/3WFCCOMA9Tbm0x99UZI7QpDma
ZEdV4wx5m8a8cwzLzi8Zr4iqDdQ7RksNEPyy+znVpHWnD8oVdMxK2MHmq/yJnGam
vHNfyzz5UP1aQiha3hloqafE8xD16oc1ion3XFTBkLn+44BHmE+rYE9ZINqFXu3e
xQJYZNEHo0AN+YeTbrOPTCkbdDM2ualrmJi+xxTjG6XvKEkYzIvMlTfOZ7YBXHiu
C3jxKrGx8nevFuzpSLTA8JpTRG4kmINCPOSYMXl4Wes2TUjTg40BrOH3kHHNld+M
GlJh5Fcx83Zsy0U6UuAwlzZZgEu41xcEZV7V7UmxEOhsECBYMBfsA1vABywiff/n
hKznENQpRRqXy5aOyW4T40KOwYTFyqtrOdDE3OJ/Ix4P/iJfCY3Zgy5fvVnts70H
PYsisET7HUbr3YiCefHSbEcN6cy12a3LpiDU4mQnqSNavB7Iadz97IlMy7FVOJ1o
3m21gB6MTYCUc4Ng45QxEPH5sRwVX8QCdBgU0wby4dyXYVp6smokguD9fEQbN+Zd
Od1zOHdKt9bsHAwx1RaYTGFT9Y0LC+c07UKGBmRLeOasJgxUCx43vxxH0rwqMahw
0wngCRzorPQO+dnjQMQHoE63PosXPTZN9oJiOl+SK5lg4Tw+qdffBVQGBhrMhx+T
yNrF0FJJU2Gs5V5uqKBhCmpi4qGGS2uwb9lNH00DelvdkbBY3hWxsjmGNersoMV0
Ycwm9fct9I0F3cT4ZCEQthOvTQkAN4glECn9g+bo/pC6VEmj5Qa4VqYfjYJj39+U
oCqddQBFvt0EoFKoP1XMu4GxB3Dpi6x020rI7bnKoKVOzwrpAOrZ29izaCEXJU/G
GoswSwbGfl9ugXPLZ/AgYKAsKjmkD7IYPaxpexp5zAbgj049HQ+WeUImcykM/sST
PKPUmzp1p6ZCSqsifFPCCe/4o+RwZyJRRGdD2LjyjDlaxLr+pwjVWAUpS/2Tx4AL
i9HXYNt6PRF8UTJsCOAHUadYx7N1aXpZlWoJKgyJauBgFhdb3nMPS4HXSCrt74GG
o3+E3IHg1RKgQkFLXAQXS3v3IeICbDv3lxa9D9B+V1k/Xbm/6UwOy2Sp1o+Mc4lO
bPQMmFWFcXBMWa43vH8Z7VHFU6MHsZUyVanZbNTOkv+Brsbzg/i1ritgl5W7/yDe
TxRaEjywh49hiYYG77225vT18n+Td78OmwtsPnyay/5t+p1it3MJhei4cjl4noHE
ILe7A2XLMrBcIklI/rUs90ozQVg3+YL+3DE819SiWOpDm/oiobDpW7pGBkCUYsFM
LZDGImV6XrYaGOK4IegCfTmZCrDDto0EM0x4PGL+Aq5FRfpvXWE7WIsuEuu565nu
aQcV/xrut5q92zPItsOqCG9D2GUUI4Ak/7lG5lxC41ypLbA/RhSVqjViuWzMklbw
JuPbCe0nqv/k7E4yWk3UHj3zJoiLlvi7x5ALxCSqu469Ik8+ZThq0iqotdceP853
pATa07AaJZxb8ElYd9V4W1UKsC7iWhsiW9hwAK6LqvEA2t5hj+yGc4PuB+0WJqqf
z0yUM1Wv5Qj13ZEAgpy0rI3cXtRR2CMPQ2coySaYqN+uraTRZaGXVuW3uPAGiuQH
NCa6n5eijsgS2UWi/KYwkyLzRQr795qQvj191S+/IGME4+sZUeHR5vqPw2qEiRQL
c3gqSsWw9hRO8tbo3RvMNpocGvpkWWZbFPjz4u5Fvsczap5RQVS+eVRH6TWCPn6z
37XHOgRjQVrWhDE3nXcH6BGo1ykcZnlZIIprXyxb2hby6KTMBwDWkzvknLkBa9kI
VYgLkpexquMGFPfx0UJCQuLGkk8PfLGknUnKLRDV5lUjVhjIuTvKK2lAoo0jHYL/
V0RS6w011VY22YsYj+xpP4q9BhV5MquOdXf5Z8rp//S1VFXJgL9iJ2q4APSqw/fW
B9aXTnvIna9b5zXpEivC1M9CjGlUJ4AixkPPWs2TiWyJIHrkYKufA7GdejaPYU3t
haXwBmdh7f0dVIIhSKMU36F/RByz2A4SV29c+U3abEZYJuv6MR7FWUQQI8JDmGk4
q35Mhc+gR13Iux8b8mrv84qbVEdYBaaRe2D930T/UeMRYLmAoOOYBjg4EyZ9GtF5
JABrxy9TouHyaVgRkeoOT0GzHSMC5GgrQuhfRFgIqqXjPswuGm25E4kHLnM3IRkj
JOZ/jQrwCdD99NaOgnDVIsnRaWzd/X8nhoxmQHo4J+8ZKhtHumXAfhH6qu6uMxHY
qDyfY5jT1G+wXMt0MF34YxrbpwyWWnj9u5HjUiKF18B//egOAvFvBZvScsF1UGiR
bDsLUYk8YFGw632C1gr1NLtIocFpzJYmJHnBPn/pTPwowKhHhD1LIt6TU5iryXuI
9QJwN5tFxsNnB6oo2lxZjfum3Qr+fHZt2THP8jq8he1vZ87/Ng9Rcng+RdTZJoey
Wcq24Gb8B18hYklq0cZCh8m05LmVWa0LJVqbogSSdgXvHmmfCAWneVsQDqI9u7ck
sgUuxoSUxG74ccLsA9Mh8cb+oXo/ygPqp3Mng1ks8S+TRDZiWjCfRzKbLh2Ev6+/
dnHULES031DUxyhpBo9wMS+NxLRyMVohZsSxYlnoAMZA43XkLdGqTWkn+4R+TyiF
gFoL3kc2FjNF7nQqnuRMtbFw+UXE1yhuWs9+yWhvQXFcH3ir0GQxF4HGY3yHgN8v
nM6EmYHju28rpJX1PTQoRBifvC4mzOS3F3A7ksbOcF/S+c3awLrCj3OIUf2nDnK6
x163E7hb2sQ7x67HNGHhqV77Sp5g5bFNJOikWPJYsAMFOu3Xncg7peSuk4WP2SHI
X8kF0SYlJE9P8fvBBAj7J9oJLqngFM63pZLu/dv2UfdOk43x82Ajc7mOgKmlxQa8
ejXp++SX4N28Q+7HBQ/6ee3t7JjyxV2oVMc5S6P3grMD38FFgTH5bGkEUiqHvYq7
OS4HTIzjesL528tJR+yXm2VPvfOmZJEaa96KryyKko3y5O5ER0v+6V/vFvoV1PZ1
YXOXl3ZopySpGjv47NBwkU/4tqegKnziPFNF7+lbpb/TpLtZYKVVi+2tPW3pEfom
h7zRFtcL/ZV7zzwzovtvsM7Rx8kcY0ecoF82W3aSAn9lTz2juPk5w2MS8j+uLUkp
zSHbhV8drAhxsctSb+SNut3K3T54vWBRjaB+mUeO4YvufpM3maUuWMC4c+tej2bi
41pYf0KrS2GISaADzAZ4QBvt8I0hHksrSwze+wOwJaIaSj91YeELjVdDlIL4HeCf
L0wkb9MGZC62//Bt5i29y4nDj53J0ZKyI9uXPGJQyjtcXAOuYuae2ANeeWvg9Rh0
z+3pJjgMXlr/DKqrQ3lEN3gBDwuWt1JDJT2CHg6faKb0GCrfM+qaa8LR8MXSkXzS
5i+Mqsro1jjVMudLEYUmaIi0FC81Yweri8xIXM8yAEzKtLnoBLZiXHA7sQmn8hnK
yQ7Kx4M63BeE4+HO08Zb/6vW59G5TiEarMqLF9lG887sHvYwaE2o3H69wOuFeL62
lGKSOl2U7m3mJIbOk9LzCN6Ttf4wE75Tr+b2AZzqL5Na2Ke4OYF0jfsc+upx/516
+mib1fVcomB25n7JwW3ntPne6q+8OnXt04cHmFuHiRUyingGJ6DZSvhUXslgIwIS
1wnw43bITHizh9flGliqT4QFSPvFQyovvhRjL1TNcP2qZ4PeWg24Wbt6nSymAQW8
Q0LoEoEYNrcwb/iqqNvink78mLnRBCRvwpqZLUJ4bi7eYFXi+cvGUdPWnDBTaJOf
mg5GxeqDPvLmd3UQHbz1g/Qldo8LwhUdltzYdCGYGgjw2KdKHpPsVj6B8825XZDt
cj5IcbyF0sCaT9CKGCUM+Vu89Ak+hfgVwdk0Dx35ycEd8WlR6AsC5oImWqRA77iL
YfzsQTcOtQ5k+v18AZSzGT6mSzkNoK0rG6Ft+HBJ/aizyT8U+nnydxJf3io66mbS
9lenNs07hhtr9XoD7CnTcuksRl2XoPvql6q45zgP4dOpLV6uXtPZ3QNn/KwqFKQe
lcgtNm0gVAhMrHPJItYLCrP6cM3B5fjH2eMSKkqgCpREqMICDUAdOmFYg9fUCTf8
0VU3ZcBQwmsOd07X8yTx53TIrfiU3LshM0I079TwPlyH2iFRkCxOiXrd2Yc9l3DN
LJFhlNemWOhaW8MXYccybSIktmn0VVUMnIm6MBerrXV5D2lG9mQK7c1gnW+BMPzs
AORyPqkiYsU1zYqOO+pJHn+VM5aN/PH9vZUmg/VJh+wbZh/EZhm//HXwRiyavBCc
9HjyhOQNWAgEA90/RulQ+Ol6BtD3X97rLc8TOs2p+abM7tMTHnkv/3SMi7ITGgCB
VYc0lESWWQjO1+ewO+OALvHsWBbbJnVDeXKnbVvu6LsSOTMdofIH507A3zLJo4iW
Aoqw1weFG6fs95tRDsDAnHI66Vr40Pqbb+YSMx1ESAWfXz0KF5P4CTBKHd+O/kSU
wc455cav1Bu6HshqZRD31C+Ur+dh7tgZCFO3EvbLwAollmcEh4K1QtYOz4xDNILW
flagF9l/4aJbJ+rD1VRfocL11j2iwJb4CiHi8BN4hdsl0XgJX+5eBq1vgNfFiIbT
AuKlWzB68f7kOZb85qGL07mrdB79qOoHOBpUEqtD8k2CUF3Aua7HiaMdoo2o22rK
xa3D9leiLPnxF+ApyCcovEL1RiisWmfqR1mQvu0sSg5tt3oNyP8tjJHV1p5k4p8Z
j+aBZxp/ELJV1iUImP6oySk8LjYRelpf1AySnemEt6XsrOAZer9Awpvu0hC2cgQi
fUQXnNoN1cLPTvzRF0E+T0VWyALIERXh5HwSHPtdCmtntf8fjcH8NhnPHHKt4gja
uHMiN4/CAcLdikhK9IB+2ffjqcfn+00Mw4zflfqIVCtbSKV/K4Eqr8MaSJ/JOT/c
qhtKRUEMDDj778EbNY7goC6uPUR3P0ZQ6KFsWyB2m++QW+faOiKMqpEY25AYoYjB
sy9svguJqPZTA8ILf32U5WVZyLQRNxs0bMJzrG9DyJeIHh+0dd1tTYXyzzAeCmWS
A2Dl7UGzwxzk4FfMEJnLC36qtRIe0WjcK1yJVTojifpbreIe0mLNrtjRuOmI/6A5
D1JSvgrteAs0L6sXfjAaBfRpCX0Ndl/ifg7ACl3VaHLdP+TXC9HOyeUqq6DRiHVo
bCc47ufwc5dQ67DaZZsSRdBT18yOK2+3f3qcSb/XGg/PXk1PWmO9MaO7PNPL3hrj
V9zi46nwkgosM7NMpVeMvYzS6hJD6U9Ysl8lGFSo3X8uYLNFHEzdUrNVUDpt/0jT
fvs4RiqssTQ/PF+1uEWJUGV8RSDLdRq2oSBJACyJVTBWyjKEBiVFkfDeQRLQpRua
VSWT3DkuOJvWr8bqOHRVJsHtbU8Xir1h+zf1IU1sIlcj7r6KWZcca3AlSzaGzquY
8Mew5mdKL5A/LC41lR9oFYhopmPgChcmQ/WPYqJf3wnqf89WYOcqGgvYkM58WBg3
D/q/3AwjQ8BaREH4onqtQ9sSFNZmwL+k/Z6/4gVgDsgxqXQ9UNlBMctu+evgzf3i
9Lq4sb0Pe17SP5Ztv91cDX3KqHOHfKr2A5Km9/H6DY9QpqocSMSesagJX8aTc2yv
erdlkAhdsNlhmzIhty/7/HC417cEsZl4giGtjk3RfFtVvID6P+NBscD+t8Movshh
7gmFtxer9fkGPA8F2BnVaCsw6A3MUyun4MMz5FsjYrlOr7683Eh0m6SnvzdqUgdi
QRmS/V73gYL4eWzLfsr3n8NE6TnFMsoWyAfk4Ac9+lBpWCJZ5r8gyNvuFpq0F4Yp
57L/AOL8piJRa8nmvc/nAncukg80Eojn1O4ENV4BABM9jqAN4CUP01vmTNUdRPek
bnRoWdTgzjzXbIpgkPhh9JNe6QilGE3lVZB2PWzvwFSwqI8NS1bHWrLNSID3/+uj
35CugoZXIsDpeqs98WOn4/RNep+wcJ+CJOi/8+7NDGZNMxbjfhZGuDR9NAo2pIad
0xVBwwI6mqryjt9pApIU+6DKSKdHuRceNA9Toyf4xeP6rZkuqyZZsCu0xuPLutRe
h83+vCPANTsTfJU7iVZLb1yPpcbAkOOJYSbIcheOex0Om9z6Bq1VpVNBneNdYk4A
RSSbyPT3g07zXP5YntKBiLX7WyZUhEaWOUi0yfqZKGknEn97viYZ8fA6YiZyYisK
ceFJcYKxpwpJQGNthFJ50e6XVSGPirTVZiupqYgfsvuFZv91Jgxstyy3qBVoEU47
JafN3EM7RSSqRHfD5gU8yryfZdLF6v/H96EGK/Ct6MP1Sznq6FQsEkvlrFsWUua+
fWnK2DJxe+GtrNelcXo5ffs4VWX0geWY1vbSP+i/1dVfRCH5YDjR8G+mk5b38ZWB
Sdma34epCMA/9+o3KeZxSwJZkO8avRNhCUiTvoODL25VZEoesdQpUh+psdRXjBFw
D9wO1lBRkP2Ufau9n78/ccU+hofbQlszk50rqro1alsUCF50feXr56Hl4ZOlBqAA
Fit2qfS0tDryvp9WK6KX3Q0nn46RAMJEdeQEBijugfcT3mMHrjVISmNK9IWL0SiJ
QESToLaAlKxs3kEdPb/rGK9vG9ek5Jfp/1jkRst9AN6GoVR3M/JY6KdEGwa2ZM47
cGu0YINXh/a4j0sz5MZge3oTNbUqRX1RcsGuQyAWe6mJonWgU3H7GVbzxhTLcgVu
mD6fKcFRXlHc9SHw15cqDEIePT3WxsNS1Rgxcp5nC51LoUxkPNilwWI5jjblGzno
bbwLKPcEOcqDE339Rn9YiU9L4TukXXW2imh9YlqZqlvBHDRGfARnu33pC2cRtL0Y
W0LTymdtf/xY+X3EZKLxPuDDiE/WfEZ1AbSQuK+WiXPWWsRwI9UOcATruUk0qYEG
2fU0UDKhs8NlFnfod6AUR+HpnjZSoIUJW/SWFzHWuyllzrqmSkPPF7vx0YxNmgk9
u/M6gOphYP/X1IsgeHgda6kYWH+cBgJ8X+onfJUmaBzEF2kqDc1ntxpFpn08H9Ws
fPClnsGv6Odnc4s58/gMneNJoeJnqkorOPXd0V0tTx1Zn6cFHYg/e6diEgJQP72E
is1Vzpk+rRLCeu6vUou2M3sVuM33knyg2dcwZbiOArS60gFX2vrUVrKfQrDN0C8b
3gnsdD+1P1aU2bE+/YIJNgdZl5DelefPGvTP1Vo1PCCjhQ69EYljxXeKMemmVtDS
ac4bCK2xUmI8bSrOC2QqxSbU3XC1zeFlriTBWVxRDZ6b5utxF4mPIzw7wdLCuDWa
tFbIqL9qhsxpZhcxjMxOm5k+n8e/vnODGOz2XfurTEmZMDhs58OCgUFP0NFzXj1e
EM0SwLhZ2tvr3fuDJD9S4vuEcxvZwoWexTZaD7LwrFjOhEo7soKm2k5nOIc0q4XR
skfJH3WekcxBenUdZRHsVqtw4csRaaptWJ1DeD8QfG6vkXKv9+yuZtoGCWmWN5D1
8PB4Pm+YXF7chOCmXDrR1TJ1jIVwFi0X6s+0E4KIX9o9XFh7fatRFth+HLANtdPy
EmzZLz9nUUsJNJMzR+Wd4lkt1doXw8Xl+FW8dLqv18hNw6xTz5a4Swxuh4FAWMtk
TV31Z8dS7XAOVSlbaLIvYCcW3M/LwJP7Mq9Fr2UW4pNlkd2TwmzqUGx0l23cERum
ZpSNy1smg8syEQGcv2XUX06GfXAzNn8d2K7v8Dv0QrVTu3OhqdN/McEBVZ5871r0
9DZNX020M8RfIx8G6yAaWUec6NQh1uj1pil4fP7Qh1Cvh+6YnBB2Y3yeqC99mWGj
+5zmfMEEC7pZuyoB0wGYGdhLz59NVn8LyE5lfmGUD02j8dQ2cmC6Tp0v6m/yOg3p
1RTIYDarUV3V9NCI/zhutWKfQLMdPworo1BXePYxIL4YzI9Xq4hSLyPmRapIPOqW
kFFC4QopjLqYru3+QB6YlMfEdBBEgCnSq1wLiwemwPdN6pQmgZydjtxoXO5TCLVI
0/99kIvfljlxBnoLRWJsoSUIZWBdIQkYAAnONTboH3/4W/GRfpQIh1GrBgV9EcDB
ipvaemu/FwDHYqOj/3elK1chwlwUhcgStADxM5VLAgKQVRUPWxswwzigptlcj4rf
TMQG3DtxVXFDKSiL1h0xA9qu0U00r+UyX4FRAse3o5Kk7n80bCC8wtaLONMBJ9dr
FE5mul/sOb+rVLRYinZa+qe9QFXVk8Zjc5NAwAoPICdqUGmVY8e0ioa4Fp4d9OjU
N2bEj3bxcZZkrmoyt06tiiDC/UNQQk8/g6wn1qlFUB7Xko3qD0lhzrDNoAA6ntnX
KpVYjdyoeS8yp2zJPEVAJ8/Pl9ZuhJ8M2jJURkkwIZYJM2JQQ0nEwmc6M0dGfhWu
YLFDUvpj+cM7tFCBsxtivz60exP3rk7VMu80sOKLOkSg1JGqMurA2AEk8F0xdTBv
7AH88er06kl7iIvaG9aT67AVpW3a7iIKfxGyKZ0Ub6OoEzaPl+foD6WsSUfHf0bJ
KstcrHb6R5nh5VfWaHIzYNsWxE4TPMxkLtfDx/z8ID8YG96yF/a3i9R5M4rgVO44
cnMNfQH09F4tXigytcPEKG6OTjjQMimZNUiG7cx8NhlmU5QoJFmFQifmXISJFsW7
zecNK2ROloGVvdMqpjzjPvaIGh7TNEtxmpM4RuopW9VxE6QMM+VFvIOi2euM7VuC
erobj2o4P5JGmYmMQwm/eDXzR4iJDrkST9OCqowr/YRRUiWBeIVq/CFMKkqRKPMZ
ygywnLIiYt705WcSs1r6+YX5KbvBKvCeVGa5DJefiyOuqWAzwYKOp+Hrsf7Sj4mg
gVs28kzrg/4vbxGGcwvjeP8fkpZ4ngnJ1cfwm8lIXsXbrwqyDxBTuhTknOqMnoYa
UKucV9CpkCq3L13fLaDibTOzRdM0lvHl/EbHeRt8AFYyUKN0uR3wvCD81sV8C4Mb
mmDTl70CZb4ZOi6JaRcSDc/VPrg5DADzN3sLmXX4l11XWYCMXwJRZOZ6XnJrJX27
Mi7dCa4oG2+pU/55coIMPIO6N9V3U10JExaqXImqaUY0ug90TIx/H9WFkiB1sZxm
JT6/4VhIFGxdoeZb4+hj2tVXKcwf/RUbeG2ZWUoMAl/8vgo6J+6X+HGxnDvnW8Pa
WBbsr0KeshwRvVJPpIWvEiqJUlfQ6g8IY3p24ICWTiwmcrxnK2On767O6y9ZIafB
`pragma protect end_protected
