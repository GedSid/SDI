// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:36 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IlJX3mq2DaueFZBUBvSG9VOsCha3TMoOROCDzPveT/826tUo+tgS4VZKBCv9sf46
Y0oI9l7kN/Yw12FjbDMRZUj8gWbJ7Xv/hZFjHDnipsCF9XCM8md+h87OapeA2qJM
BI7rm8mTZdrtVS7Im57HgUndyPzucITKOCqshsMkd60=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8416)
AUxRfzWHQlRciC8KS3rCxJ/mqLj9sGyWs5ljT7KRgkJYbJlbGZcfFPcthjChxPBy
sChPctp30GjL/zZtOwne7M5VbgD4LOdqjKYmplCo3Da5QAWOXNnI37oHv7UY1P2p
nwpfGwgalNBKTS7xWnks2Diel6xDaoqU8Wk6WraT6ziaiSQq1eNpQOYBISl2B6ZW
klPT/wWfYsdtIr8zUeOfMIuDKmhp0vCqjTxsLKfbCsvdW2k6YEu81sd+sRCX5RLY
eZLNeKRXZ5cMtGjw3Gqcp/YLBVmuzBCy9vgY5SsGOn5sb2JoRIBxNUfOhKv2f0OL
76nsL1B0/EGs4oL0rqZz/oPVagLiO3Pe9ljoEHLEt7IJN7pE/vmpPHQtwZr5XTTc
01ukdnDme3CiczkZJ/KKdLCrkeUMlvu1GFmTdT329GICjQyRMDhOM0dah4LwKUzW
IWnJn7KtFWKEVyFMp7sCV3zW62MzhHZuaELGiwEl63k8ayU5iFMhIl33ZA6fFNPP
7UrfrG+nf8fSELZTywgFp0HtRfzpEmaxTuefvIVK5YkuhgzU3jXqwa9SNWsfXn8h
DDsjrEDWfuPtAj/4fBB9lao5A1gQ99xmPkB7yI9OGsFunXYNJGX859LxNSLV3dop
UMIomaoq1hC+GpfYWW8eATh7uyjmA0GSynzcOSbtfVSNk3NU2p8Z9xok2sNrFvAi
6i+c4SwPYhtA04AFSjYRdwrtfq7p5qRJgwbt8UKMqijeyCSf5liuL3Q8eBfKimj5
kak6A/2qhGl8Tu+6WcwVWoIoea5Q4f3mEvWCvgMNdUzy7N4ab5aOFzl70F0FQPdH
EnQwHJ8fox4Ngf223h38Apl9uPnjdbvNNDrg8Ycqe4zUcoaKKqpXatOcwuue/zED
HifOUyR8Gk3AgpPA/W8ZvIY/opTY+s17j7hegakmd/kT+1zouz9GsLROiBN4xCJK
+yGrLfo1TqMAroHYrGvQn9NfcgOkBQCt4oejvcb16002qTJ9VA5WcCkHROOjJnl8
JYrcHt3B5hCVgB6C+HbsFVQi+wDw07ZIY9bHjt7L+jMMQ7b6v2+QhYm6LvU+YBuR
Gr1Qec6wPi8eFYWfGzLS8F+F9yKbWZxy6bq4LLXdDNJxH1bRRm5nLpXTQM5GCH1G
joaWgwMAOd87++Qi9AL+56BYWDtUbWC/69HAtGNSrlCSxDi8UeNvme4nVPRVcvXF
+WIbaEsLj8zTMywxDUsH+y9tDYHMxPBLSu3sSgH3HcY7NMB32pItq4lLe5j1cPSN
a/X26gpbRjDPjvug3+dT8Bn0k2SYGLZYefkllPWLFYJC7y+LSldtOWSiT3V5JUS/
F2O4IVdyjPBEN1jfEj6NlbZvhvH5sW1IekSxQDyPDrULkY32hrGCC1V6Nnu9veZx
hIE3FCQ/n+VJJ3K3smLCsbEXHww/mOhU93e0Z3p4G0DPX0jvWuc5Mf1Sg/fCUyyX
3qIhi4oEQTQKvrMK1KeHgR+VNkjtRFWvWQfDkkWi+kgTt/kONJwV40HqsWCNeQD6
YvVCnNDr7dIEao7c68gDowNZch1OoH+4Sn5NjcMz6+1ErZNjOCiz+UcAcf7vo8Qf
n30EUzdlXlbO2QG+o6FIq0yQWTxdmeM1LSpOMqL1Wx5ujlbc8+t06HqAnzpNODzT
SykSMpEHrMcXBaLxfvqxhfljSoJOz2DPlPiy6WuLPFzhxusMN/yCTf6P7RV89mX2
ZEkIBL8SqrHSFSjDWYRnsyY0XzjHvn3g5U2X0FrMrRe06nKo9nMH290ZdMvm0sSs
m6b6befbp89IFTkK77XdkjbL5jaHnL0IkTwy4ufpTtMi/3wg4mWf8TBtP/iumeb8
Lc8MY87VSQwF8f7vZDFitbgZZr3N1CFEnzljt39P3hUSX9qcdVUiGnw4+f4383Gp
WuDq2Jw3isOD53T+DKyvVQsga4MMidsnVnUWVKD5eHl1UIF5sUw7XxT5KbbIqS2g
uYdpmNgIff9IW+4hgyqHjJzei1yC7VUJM+doakUxskuHFV7EAsXd8CYmHRCj1JcR
ZEOUbs03uHsF6QrTiVnoxGi33dfa+XyB7qOwuyhaUCGEvbuapGiFWhFyq2JPTFRT
TwpVfKwSXS1Dbno2WK67VzbKyKXS7iHhHyZs8pwkRH1jL46mvjizHyuOYfmsV6DC
qVBepuamJTAvw99WtSuPQF9rjCuA5qi9krM6dZeH/30IrjgAQdWCBErrGNcbrvc/
gIr0IrHDDLzFYH+0NDSoLU6gyreQnrMP3R3iLv70bEhK2+byBZ7zB1GCPU+nx8H1
fwdPXSIiCWdo+uy0QBNIFlkjyoHiTq7xB6VM7JOOd/CMnBrq7owQ5EW4KlWWlMek
+8DSyKlgYvYClbnZcHa5jOlCYSZRx11QTifKsVSL+p/cmyEr3gTM24tjT5fZM8r4
wVFcbqatjcWbrsd6Y9lxh9gDJGU68GxLDcsC3aZ6nkY0mPktHd0K7S0RzhWa4W4D
JJ34+kqCfHS9J865lVujQpKFZB2QyvbPDO+A+tG2I1l1ZKCPegYXK1lrzzk58aqV
o7J/WDb75pmbtEI10YtgZzOA4itjKw9JbCSoLxKeVg60embSGdiZaNN/bD4F0u1E
TzTVcMBSAZkH2kLUMuFaLvqzT0Ds8BJJebxx2WDeuBvFVlM3JwgUKGEJThz0XVlL
MB80eKhmTbiTNFZtW/uedduH3QC57v9XjdxLkOH3FL8qVKzbG3/ZarAu2q2kCBOW
f7FZxR+aXQeYW4EVf4QUpJHtapq9uHZU8ExIB32zrsyRu9klnXNylwEyyVMBI9Ef
KR1g+EW3fbMCRBUR9qddTTIHGVM7Jp5Lec/Iu5V5Fr82mEQFrGbD+mE1D/W0/Se6
0e8eDsxl1W/2mHn8SoDZcyMJVTYjQFdbMwZkAcvCC1bOOEvUS8OoYocrn2g3NF+L
KtoyDLwDrYRRgsw5ffwCg8vWMOBgRL4vTa8z8MsSeWnRY2o3vkEozcCY2XX6HgqN
/FMJJXPzZEWLV9PqjY5AFwmrtDyQJDdyFCYNI83DK2wn9tjUiS1L49TOdbEDWdXr
TqI0PW9vprDr8wSiG+sSpeNWYCmD5c8e012zHCQYaTY/gYxJKY9v7grD8l5TCwIC
EGa3ynFDR9X4VgJ2zdfjvbdj06QJKdryvZrcqOjFPVFNQqnMpjU9iTu7vurA173K
a2Si/7A9LGB5S5epCnA/6pWCZ54C32j2KU6bAaKLaUCjLl+V61CI3/9KZpOB3mim
ZQ1vI5XFqyZ0sgLKye9emuvzIcfUlhzqNwB/0VSDkDYxpo0ofrqKXHJDSandoJTL
aWw9SM7HjfDUF+vJ7VZQvagTyb6A3MXr8QeN5Aul+E/r7azMP2X0GrNbFlH5eAxF
D4pWs5sb/QVCzARRHbDAajL6WVsqTZylnfSI34WwUjdEz0gI23+78wyrW8GzzAf8
GmUJ0Bw+WntQH94EW1HRIYWY0+dZIMUgtpXidxFpmnSu1Ed88rM7HjYsOdkQiJn1
xiI7a4foonZ10BW323zEiLfUjdcE5TJXxh9qKBK/Lb8Zg3QHrADuwFlhk/w9EI8z
6mzO1cUWagRgiJxR9+Hr0gf0mpwQtyz4U4u/mkl7pjkyeFXqxQyD7WOSr5fNZQ3a
4cWlyf66DyBsCKrEIus503Tl+Ne+0c0OFFYHUWDT4KtZrJNb33y25Zsec9c/K8xg
KaOm09L8gIM8/VKwkj5UEsvQAkKN/GlZ5fnFUK3TnBGMSxqQZ8D39UjnLxY7+SkY
BnvKCGL2f5Qq+L1TViqG5IWuchHVVDVNj4y8dT+Xtr9AqekxynRjdTmU2umTVLVY
4iIhEtAen3r6B6g91hNNpw8TXyquIIOni+NvVQ1omS1gX1jmVF0h79kLgVGmfHvK
9c04xaXhw8KPE/jSoyR8uDzxJOrqJtVZTaY7yasZiA8h23MsEUA1CpaK2O6O9tce
BNb6ltsVpG3yuElTcDM+lKRbfIIpQ+Ow2qB3oNHX0ZaqR5NxiPdJ4L7GG5AGVxPx
4Isba403wpVjNMdjL99qeu9o8Ua90Xt5swaTcEfm+PRMt3Q1uwl7gbp0LleoXygy
qFUSfbUfZ1RFQS6lRWfuNFMKAqmA/4IBVZCXxTDBXFQyJWCzav3a/f4SbRr8hwya
+5hfPJhW4HgBx03m2DpB5MbMQn5MVymUBqZdZMlTPSIU2V4F/soIdGG/UoeHqBCw
n2SyZFzIFCISg1MdTbGCY6yDi7fmkiNdr/9uPYoGY3xiy3+ljIceYovSQSA1OOVx
FJoiCKC28t4irgnSfbNBI4ZIwxhxM/S7YYzFp3HxuV3HJIL2DxM+ljAiI6YfR44y
gtjweqbJ0G4YNcrYRn/tLTb0pVvKuzP5Z5nWmKxUzsjFKKcavDrtH52pHl2z/hap
3xeOwCoOyoIJuNFWqmwccDrVbWCsZdO0HG5ywjbhJeBdikNWN82awuH7NG0Y+2tt
2VfdIn6jDlLVMo1+TAyZhBkyXoQ75e8GVb53R7xSYQVImmdEvefjRu6UrapgRDe3
+RmXIdHd5W6lciVyaGkPfElDhBvF6/EDEBr59p8HWTlIb2iAl5lh629UlyxINZ7e
VZikbMnDeMBnVrMXuktfdgKStxoHctxbRG/fCtHXgAH2xdOB594BFQuI57i7QMk5
xctyoVjSbGrfO/0YWn2+6hV5BLcV58mS25yoAO1Lz1bJvyJoixisAv34A67cDHXz
ktyRGuF/6DJDOBnyk6p9TadlXzR0fYLB+NFr7B9o3ZJ4VWKhVGaMV1nO1uzZNguU
3rHfF94FHth6pzePyD8nfoVCNE+GINwAv1vDTqpVPKTXMzaQj8IogFdlhtnr2PEh
Pf3hDjQUNJw32dvZGP6EYKMElDPDN2pZVzhhFHMvk1XgKWtu+5HRgI+A5O9MT/Yh
Le6AUoHkxYsWEImla+iJf7kLN+hL6RZ9VEOFda2zq/OPx4hGjocdUSJ1qUvcJuzN
lhNV/oIYC1Bop2X5HMy0J+eamwC6TF1PT9xlfHhX+blO//o0g1wCwJd0eqso7gzk
ywS9Y1ywtCJTJd3NKrNpiQJ+NZS8VcyCc7JM+MWT20i8a9maQSjObvMOufV3cAXq
Z7uKFPjE/kM7bVd5ZJgc12/0prJyMYY8YH/Tjubjw8a0aJfLMaFPpNgRTlZA+evD
s+ZKIbArwCnpL52TQ4fezh00j37mawY6WYDfpRLnBscrGj9zRjqlEix8kdwWeo1f
3FeDOU82KuwJKR/dt6QzPIFMEAcTCZ8mdRI6IqjrRtWUexuPliPq6RI3D+qIU4R/
+OldQY7gZshkEoFM/lTQGvB2fA//JBbPsMaZvS6X3xHQgC1t3vZwfYtMFQr32ya9
hIVE6g4CRL9agTpsgiuMhgEV3OiuHJKVzreQIQMx9oEVcKATgJmdaQzfH8sUfPKx
sJ2TBNPMLvjdoskwH1nTtM+TfZnPZD0gKfaocBtzlZAu+h13GmSnQxxc8NPGpHO7
x6IeQJNYjvE4Q4VsHf5df5uy1/Hribsb8C5ilB3iEe/D6wdQL/nXG2ir2S5vXNpR
gSGCcJo19BREi02i10VXHo0Apbf/VTEL7xlGw4FBDpVHM1/C41lt8HALOMjb/A6+
l23K+43wdv4l3hp6yGZFjKyY5QLe8VkMEY2w54ULAbUzUNNPaMpnH7qaJ8izc5vI
iIXWC5D2vybtCVDxPuIIZ2Z1oSUfMEMrCnWmBFqPV+wheyHg/71PNFw3onpidsId
ZJLsDwvUOfSYmmFaFOUYnUcVBf6N3QpUh0lJfL1qZdj/Ds44naiSYElTK4SuHw2j
F81s8ZxEQh/R9YyezlCN6xS+YGjpM4D5W/SUP9uFK+p/g9niiWzyd954vWGTfiym
LYMF8rvf/Ek4Kd6ikx2mmBIFOqHb9PvobUv5++ZcR+cskfLaYY3C6PUQCO6pVCgw
8rvxWiEaqelusJSD/IimAuxpRRC1sGw5YB1+YHdyxVPzDySvRyavWdLAUl6yhJzz
8wVIHx1KaByMh9S7ZBTcKgy5N8gkFrUlI1zDB0st3ghVvx+YiX/NK9TlMVEZk++7
+bVS4In+j1YWeAYYjEQCKIvlavcQ2XZwzbI1icY4NGu6Q8ylkcIKr575qvCuof0n
JgFb9hOuthVaealvwN/zAwORlNDY9TRv/hOZqnnIfZf8R4Zqqrt3V0ssA0pB0n79
FtiOwsBJiEDPn7IxF14Z4SASdDIx649AiRx2mHdU0/JM2u6MVAPUMwQcbHiVKU8V
IzQuSu7gS/4BV2mKMKl2lFZq+X0iZHNgAxyWGkgRoiG3mK81xmaZeQaXxPqTA1sE
VgMGQAWb+wo3lmkYZUW2sFkLaz1HIXwsZr9YlhSt/3iz2/S01RegO0NzIp5uzUOc
dAEISX1yVARw4fe58RQ3RRoUbEuWRIC3+qFDZdGhQPaAV3yqZdOraLRlrUTXeePB
3HqOypN/ctgfMTEqCo1hV/PtclVfcctCwiFv6n/ihcl8kM5tiaziOD/BwBDhMsIZ
AWFpK+MHal3iORFvOLuPnkbUzdpjl78o3EORWb1vEcSb2hy6I9396HHwA+zCAXRc
UEaQtIeuaV+emAWp8PcgPVKD+7oB7SKBCVX5mlXc8yZm+f7Db0ypp2LRJ5MYBWBl
PjTTKm2wiwQJpWKXXHHHVD0iYaxNyhIuARFpyqQwxBk5yxCF8O80JTRrWPVObxmL
7FeR9/EaORE9mcQ6W8F0Ez8nz4oVOTxxAF0r3aqw0hGchaiRTdX5hQu4vptOxIMn
0gE/VsWMTdRDtDp+byGZjtFBuGiqR431sgR7PCsTIB8oad12YRHiQbgVzI0hTEcR
whrd3QF9eUZvWMpJR1XlPCIBfw+skDR7jT+kaY2DkpqbESJbZ6f1shcM3YIpNwZL
wYYIKsvFYoqTeZzEbK3E2mIx2OBj+rtPEq5v5J28tqmJNffTD06tp+8Jqrx8hD1r
q1hgbNHMC8y/F8aRksx9eXA3tUANBzjHkPFTVcNgJGC8QzKHMgYIQZIHXylH6nTJ
87doSgIZbnu38X0XElp9HQbJNTW6QhzbRtUXkDXWiVQXlR8OHNW02CyZ42oAPUG3
ADsJ552urk4G6TlcDVFoIpF8gXcgwBgRvKAgtZYAsvEGn2fdr61A/d7f38AKpmxc
jsj1uRNeRCN7bYzvQUrUhTBfHXBFI/rKxeM1b9LiIZzMatnucJBmGOiimr03SWEt
ZZZT6nujvL6q+r2BWpFL6Xud1RV4ZMgTGLEwXIiAKRtiJv6gimLHkJJC5c3KUZ8I
d8x3h0QMuYN54EDateOf81fAuA1gwav2V5DalVgOyTq3qzaQjed4o+PmqXwksNwJ
xggVKPFDr+0/YtaqXwYto4lqHCHkL6ksdU0fLyerLBPw24xxCyKPVbHrFwxcfA5f
A8CRKv0wwMeEGE4SKJ3Itv/R0AEhMhc5Qe+JnCtdupMRj+t9s1CjahhYjUM+ZH4k
igfO6jDZahtlKexv8V7DHytpoMEydlUNQjkgyNogtVXpdPM9jZ8Q/ICMD2BZXSl/
/Vhn/lkkCySZ8ewHcfQNywS1S9NTUESzJlZLIf/zct8buycZgg4ySy8KxN4tWUGU
mgpX++ouU8TVa5DPvUVoT2ZhdNCs943dM2WW+OS+TQ2S+0l4fGK2xDkRqqRX1PA/
ODwdyADnHuyEB1UihIWddPqpfhqpwuBbUB3FgY4Qwqx3ESB74wgY8+YR6lrFdo3N
gWTJdI0GKSztwAerQmuWNf/7nj9/cBDp85wz7NKWsTMU1SfsqnufcFogkN04ClHt
WdmGItWvhO0yyP5Ulo6qB6mvd71H0ysWHTzIRiFUy3z2UZbKF5GYmG+D7ZyKgKzN
AuKhPxGPTbgksziUZ5TaSXYK4ZKL2siISUKf7Wwo3r0p+/f3+Bgh6EfrdJUU0qE6
Uk0cvxtNLh9fT1N8Pg9JPWpi2S7D0i+2ftKHqVuyKnmefRBXte+hEXG9Vm5TZLLG
bllN/r2qDaOIW0J02+KooN+C0s/1eKYFpzIz/EyI/ysAeRl57QS0ntFmv0+UlxCH
BuXCvbuRrqc1egmZRcTHAaC2rCffvR2gByZ/LkFXey6/jU9bfB797SpZwi2tD5rM
xRkzzjxdxaZJWctaJxfXpqfxAgI3hHqSVsOxMGFmYIwlRm5GBjddT53gyqLEuOog
nU4wyoFxCouk/7QHBs/1GTBbUHXby35Z6gZ9Ryl0BMMEaJHCLdcmd9/+4oBSPDhq
XT9azAvCbz7Jsczl5QL4EcYaqLLoix5FKZCs2PAgpgO380OIrvCTojxTjKH+GhnD
cLDgWKziLufpjOBZYQTpK6leQKfrY7iSnPHV7s+fiWWIkWQENvlEdTzNot/jTbZ0
dxjIM60CfPnvXA0v4/Rgmv8FJst/Y9lsa7wLOTKKMVusJXtXdAHkgZlDDlPeNhlD
kH49hiRckzxt8pdmwTBFKMCYsFQqn+2ZaQNKWqTEGUc3PZX5xoHLJF0J6mGWRuMm
CyGJHS/Qi37Ms+MdOZSBZoc3c6cnyMWNFpGqdH7OggX8UcTjSDmW9/GT+20tz4ug
k6/o8u3kbzLvLLotj3D2RdL2ISgNnJUBW8s7peznfP9iGrXgUJb1Yu9MJ1tj07Ad
ISAjvuhwVbR2152PztmyXPRyNyr0HxViarqU4dBIGnv46I0Bf9uXZwLdPzUdNlMe
quznN8JXjbm0XwwUiiBj8uTXLyIpMqkbgm+pDxwNbH1IOBxb+ErTqyFgE+rBNpWo
XN2xjWgJ8ZhFyEd5ujb+BcZnfxbOMMYGV8WUo2fhPoJHK6c6bYTMqTPlEdVBA+PW
LsB23jIEFgEQS7MZpx6Z/9gwdl3SYnCAAP3RTfO9zB+cWRl2z4o3wXTE3cowtMj+
BmTpEh0sJNgLiFRlHj1MIyIqSzHKBoO2a/OSYq7tjCRMa+Hcs5qcY+TGuU9okBV3
Wz8NW4RkC+/TrSBv0LozmTya/oWIYjnTLqdcK1xHFHballqy0789o6u7396ndTsC
XEZH98BoM1faw6bw4txSQpPLbgHUk4Jg7ghD9x/kP6uw89bb3YqMtQSg9h59U3EV
M+JNBhjb0IDFmZ4NZgN2o5DxG99pOKgWUGCtbc5bYh3llwjOw6Jn+Lp/Uivk7hek
LpVOxNKPxtaS0tCZsw8KbUNMrvAUyQxCrh4w8pnSD1qjkGH7YTVsRAxxxBFU3LEs
YlR56jA85AwoiocUFkmbZzJf3wpNG8AOHSa2DkJ3HmwguuxPxgwDStIPiSMEQmaE
uUiYUN74k6QkQPel/G15d0txchiRSeOrXGPw0I4LhJmdr1MV9opGZXt+9LtkXZlN
4k+Uksab2DppmFPk+o7h2VnMJ3B2aGj5OG6DMFXqanQPl38H6g9geltoF7lKRQR1
jl6IX2nsFfYdGcZsU2qGqjKDuDzUDIynryKsmI22+kO9kBBuUpI/Vwap07E1s/RK
lIe2KckEwLUih/3wblJK4eE5SJ0hsSWGiyivuez06fPZJL0D8ccGLmGAeCbtz0DD
TRAtHbg7Gdiq7kjDsbIkhMXotKujU9wV4jvoZFo28GfsyXRQlqN7xal7HlVz7WPs
X9+gD01aBoE8JOCyNe/PL0LFod9ROH044TElLmi0nk5nAnBxflGZW1DP6l6qR4KY
POFsb/ogCoeRIEyVGVPPeTylrh8nbYl+BKEmn/RBvBinrwYzlDJn9QbS2l6vHx+W
oUqpCZUGyJttEyYhwp3xeQ88RsfEDloJfecmsL8mqlKgk/27x0ZASd8MSAMtJxec
jSv/16v2gYcfbx6x201PXn3JAyq+YxSEu1f0ZXQX9X61oY06qXxSvQobMObTa8Jc
e6ssOTA/apL5Qfaf0q96hBgc1b37AJQ9HPqktCSLrHeNiqRtnNE2JKvCVdiTuG2/
kKKVdTqz4bBK5xhyF4yGdgOM9eol99ZjraeXY7wy6tmRBoLnMg5UWBKidkz7zrPH
ma8SqIMpzUOisdqBnaYS7U5FN+LNZK0bFmAuUtAMVvD9/mXvStHYPb/V2DYpJDgT
Se9Ok3A9CAYbPoRwjh6qbkQFGJyCnsBV6KvtYLhLaV7oZ4zCEV1iyy9ZM8k4GLFx
LTWBfKWj9W3kN6Xy+W+I2q7zF0jpPNPP7vYdWwVf5hk0pvyRy/RZD1lJ6BxUNJvZ
liz7aTKAFuGHC5IbEWTxNNTfPyTzk8yL5U+tUfTjfAuSltkmATL4B69w5La7zt5I
zA/iChvDQ7us286m1Z/q6c2oM5t856yGa99MejdAl1iSlohWMQUd83gQdk8VIx9y
rcqtnPqV8Q6m2RfhPMjLcof9Sy83wwF5lter/vTw8Uo8wYMENlx2iXau8xtPfrLU
32oiwdhLtgy/wiSTVL0iABJrGBuSAoBzsRionJOvrGDGRBVMoHD/WDSboPOYIus8
qd9zwncyvUUXn+Rn3ccAkgqWRFEcqF7a+3P9sb6YdnA2v8ACH8zU11xfzbAqo8zq
m3mnRl6PAnVEhpflvBysCe7TqpzGJRBuYGKthh7XdQWJ4B9qUhqbWkzjswGEPfv9
v3OL8gOEa+C9wjucKnn1uc3e0Ls0N623vMSjhxcXoAv4DY3UYcX3TBmkKKn+ijlA
qRODr+cKBW8Jwewe3sXVadoVaHViWQhJbLLSM/+SZ0A+bwIIO1U+1qBSUV3S/26m
iS1aLnSfy9roXVYs6DERWG8k+gupUeudPDiTorNdVLGBYz3pJTXgxaKpsmhinh1z
1I7J/Kvq/fW3+MipmwX6ZNfShpb/VVbBzeGYKIifntxkaWJBr4Lc+DGyamnqFejT
u2SE9LOvouV0sdCZw5azhS4NbodxMQdTo+MswqLWIaGY2QmVNhI7CarsiV5NKAvC
jeDJnOaTh7W/50g95oSaZ69AK8qvcbJMSvx9GEN/EMMKMtgL+elEoMMQNFXG6WNR
c3GQEfq9/oYFbWXHIrY3uvI+C/KNvUGNNZIur0GOd/sWOx9AMOkmnKM6TBU1TD0v
dXCBZtC46qCZSfVeeX592Urpg6I0+6m/CQZ+t9wQUTH8YYmJ/ns1ZagFeDALR3io
02eyU34T4imEtU2uiG3lcI4P2jfBzx6M/0dmCVuhy9XuOCVZD3M/PNXJz3XRnfMr
VeZZBrINOxK1D93uUkT4QH0EVVaw3AY20Bdxt29q8V/7w+tYi8dqamjWRvQ1EFz8
pWIA5HsEsWNoOwq16MihGQ==
`pragma protect end_protected
