// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:35 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tjNDy6Dh+7TbYzo8uPUdQedcKDnWAW0xV1Iu7ax8zLrjUl6SWZxAxORfacfpclJR
4tTBfW6qvYW1bEO1mLSwWwjCOAJXVNrlvpmrvpHj6W2k2pGkZkGCLImBKGT/do7f
nfchSnDmDjSp9WP1pv3uRWQAmmAp9liphLCqW71D4OU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
LHKdvMZ5kfi15GWfJxB8ai75S0KdC0WyrVwzxci92oa0JqXJG3MgIO/ZY9JTAEEI
Q0tqC0L6Ac8Qa1b6Tkw2cEPEySeLVtK4ynGYxaOrtlc6oWikykVHEvmUzvy9V6VQ
OuC2l19lg3eIHv1PoFNzBI1yyyg4deLkfat1+PVfWce3A/DuEBTEBdk5InyaL9bU
89iMuCX2/FvCZhrq0s9MRaPPAP7N4lbVmEJi+9DhIeHxk9T+TPkjLv/QWASHdRFt
taQDcYrGIiGG6u+JQEmtrQHDt6C1boCWi9/+CvOrrbxQkjpyNz339aDrgQLGZDs7
KMJKF++//idV33DiCrtRP3iEHmYvoSpXItkqGa7wpnI/tUV1SZzi57MaPqc+SAA0
JJvAKzQSVA5c/lG/cdVIFxRowlrjKLbC/NGZDB+TarL0HBeRIDRhQ9aXXRcs6v4Q
9U9T8udIJk30Z3NP4z0tmysugA0WmW8gCHjNkzu8GrWi1rfF0nZq+wSaR1tVRx5Q
JuG2SYnufYT1xwl7jEMimhcnUgdsgQTsqlG8YacwKZ3irJwiAE+6O8EEtmYDM5uQ
4zNUfODogMdpcrFxpgTO3QxyQ7DJfeD+g1E9c4XtCSYYmJUt3WGwPGe5TCck1BtY
WM6QoqrnqO9U0Mx0tGo26F4tsa9pRqxAB0RKLiYNvXHjaX5/9BjjfIxfRXnZtjBs
c1Nl3Z2INPFo5vYLs8cFFL4PLzbljQYi3ttOeFJrS3gk/GT1mjLq14R1VTiDF++z
3ZJxFe/oaARXzdakyNVeInU3Bp1DGxrUdwr9lN1yBzCh1Xkd4a5SNdUbkmCT69KZ
PYbBEu68f7e7QlPjjLeEGXl8CUm4vBzXzkbHIip9phTlVBFhVVFEqr4Yzh9SAXYR
raru2pTT6eKMdAhta7RhJn492TjEiJblWySMvJHd8Aa2tzcpocmBBwVnwQPMZT0c
MHIcS7kkgJ6DXnb5Kt2dOVIeiDFJXzyaeogZiND36pNv8eohUeHYVJ19jQh+A3q6
WHdoZdFBs015zrtSpiWU5RgjnyxuuhA7Y8MY6y6pqjgX5hIucIfExiIj/oQnVERv
b0THmWO2SeDCwfYE/qBC3ZdJ/wvXTRUpasC6OesvDTBne4t57ReE1z5APuimwEBA
3ly6f/cKdMsE9Mkl/r/zvRhW8NIt5LKleggzHKcvBM7SZ89249yNqgRfoCzAR+5E
pXnDsbwR+M2qCvJo5ZC+5t4DTAK78cPBEcV1UEU441CwF/VvO2tfn5mmSxo5P4lL
VgsqBmqaW0A+2lYc+gEHvZ14SHhzsm0YAX/+fLf1XdwQqFm0Q3dlIqoupqRGsWeL
jgsP2ZGvbkg27DNrTSrjPaeE3RefqCYm+ulBUkQ3LBAEf6GK82e26PkcRnuFFjnN
nQrdvfrkhWw2Tcznw4kDBRIUN728H2+nRCVCkG92pR00RdsanxLTRwSU2/fT8iVV
G5VMbEdNxtMUI3IgpWkkAkBm5SoBFcwQhvCxw6ByRezfjLyA3RoP0G6PGViB09vA
Ihz4YHWOzH6pX+dS2Nx39erBcG3YcwMiopi7LLi0oM75QOJDWRqg2kJwtsZKJqYz
O7xGfUEXAzziFd72BUXgQSIihHi5BhpImVnOBkeArt/B4LZ5fxUtBOKGVhqSJ+2e
JF5hgO4v7etI0yKDPh1+oIiE2dgUsYJmLvknBjlukaks6TfQZTStwMUx05ojBBxT
5kWgqQVSnTfCfRwcnknTCKglf9iQgJoLPDuUYD5TD4SHuuBY3/SximZgETR2l/ne
GWD1LyQuvD8Y87E2Pa3dOsg7PEik/BAhq3YzQcWWzf+LyNQ22POACkwoq4N6W2jx
K8xDs2Pxj7P+5RElDStYzWw8d62lu1heScNqWFsSi7o3p3l2Ui4WnYlqFNcr014G
p0+U5ERYaD0+LTCqzAYby24H9Vi59BNyuvorWeRUbAEMQhhvzCKH+eZdHK6zEWm6
k8aEN25TJTJQQFgzlsN3ev84ypfoNgZWimMZrOuScl2KD+JDt+afBLq2gwv81sHL
U4+Ist541g5OoXNx8jYL1vZV4WDcPQYftNDGx7W5ht7k9OWts6av3OVmCLUFzxyM
wXjod9cCeg2okfH8Auk7r5PFlFY46mML5EheB885m48Ss13ATHe4noEynGK8PRnk
k8O+FYissWZ9NfVN572TdVuZLwSENncNszgdaYNS7RzlWg+Jfuxjst8ErApGKPLs
SOLnbZUWIHTaMou0t13eky0ZDPB+lh9j83YTJfu+NKdU5a/4+kX5JwRB3z01I2m1
KEw/W7WjlpxebUHYvWrZBeigDL8YMwP1kktx+FezoqpLFVg08grPhf2N6AEd9Lqb
UyXo991FkxfXma8LSVoOxIQWQL+8jSi0SEeinQeQuYJihteM6AtazquciTvjoaO5
f/lVCjO/Zp4F071INFBrfoDGYHKpoKMrr3s/+NEIcPyQKtIeo9WcoOZqazA1Ttmg
DVCw9tFeDw7NJnEPm577W1y7c59GfXJUp1BSav4FoaE14fP4CupJw8y+XnkhNdDt
YJYJ+wEgXqJQicv4QRibRYFoxViDxqCU7oLEGzc+cLMJwLhqXcawV8/b57VMD33a
47suCY4cimTq3GEBtMNkzRK2yK6L7G9BaPkm9pXVIg1JP1yC1+0jd/p2/3j3gHLH
yY486dRk/Se4rODWanwuXEtiAL+bEHMpaRMHEmzzmE6C8499L1GHKWM/VG1bj/4Q
T3f4b3xsDUpynLpBUPtbpqkyhP24AwggUT1Ebs5XEFSs5ucVKk2qToR4BQAXFGSS
L2sX1CqfQhR/5K8bClZt3/lhXnpEdpDt8oCDYcpVhaduQewD1WQSEDAgBFwjjudj
zUuRs1waqBpJUqhsi62KPd8/kfaEX029T8ZvQmW1RbBD+f74ujPBpOtuvBV4m8uH
35xuz7pQIp7UuuhJAZw/5lKuF0t6Mx59M/XQWJG5zqC+z58hzyQHgUoQsgX8274M
ApEc5ejpRUgMrRgW7r+z0oAr+CE1qis4XZDxhPu2pX0pwxGn567rxMrQa9fZhm3E
VsJ/bU3smQ8JdcYbZrEBnCPKJ+KpdXspsfDIRd6QpyezWwz+Mt5r969hmpHH2/dc
sZ6GauFNbvfGJIy7h7raFhefUDqxRLIvtto7jzeY104RjC4vNf1fC18q+4lRxzal
X19OSEl0oum5QVtDcUrd6NZ5mPElcWqXS724jRTEdEQ0+lISkOWMhHf5iXkaIq38
veRke4USxGRcnEAOETy+Drel4937fUsnFklg3QofZxfBsu9+D7ULvVLcY0tLQa3Z
oXCgYTWQlnUL6jf4SCEXAmzMMnfhcYTSs7h18Y7foL6/S0FBQmvmeoNIm458D5if
NuU1Hp8Xuif9lHrVxjeD215HDfDcjyw7Ai52Jj1YZwYpKWojC8FIIf5/WyxcY8UR
dKSPjUSSvEUY6eYjwym7HpM83icPo4SWBv3He44V1MpkGoAmLFPk9WIdZJ/ltdFu
kOnVtnHEwnsKxImygCGz8DDJGLnFw/ipCzouGGx3cJKdO6j1WAa+AoXV+MeponmS
pA1r2TEOV4NfZkMDRha9z0dpUUqVUIjqyHkUEZkjGjMuzww8eU26gGU47dUm2wjc
hUupYeprJ4GWrSUZpBPLj1hPqM2WEgQs7JIKkeIckb0ASITKi7x6MJnue8F33er8
7KvfbdBrgengokB5/JqalSCxi0Tw5OzDElwejfiXajAfIhjnZutKwZVPl1XhUWLV
uMBkqDjvo2rcSv/ggh39hr8lbbUi2N4tO2wSIUeAJHYoX0fxTjcMNd7OF/OOU2oD
c9Qe/jLij7Uh7vbkmsosOGRQTTnCPRAesIBK5BDAWlW3sYLa9aUIrM4YqJlickgS
7EiD1eSjQwCpYGsD3wL1WvGXTkPSzaqnSLfFo9g4kUPQjeUKbPF+VqcvgdLKTTaR
2s7n6imRdiAcbCzgwQy07EHqbtICmIv/RdFKXav9TmZ6nnHIgfod7ur+EYDPCyIY
aSX/GsYXHZVYvMPIyi8Ol203ay6oEO849k7mGdnftGbLpRbk0CIkjxBOmZzhUwDH
TRJAGu8mlbRTTrOgndNcoXMepyb7w+cjjL9EatpjZrCQCUWiENWhuk3+Dn528drY
GljKbJe76PV5ubs3vBpa0mlOLbrO1/kykFKc9hSSnfkcgn0LblGnPtKA5/Ac1e/z
tNPDFMyjzFgvskzpTQtbHSuhPAtlbNKQWm6+L5aZXKS4/VP5gY5nTDMkiCvUl/OP
c+7Ii+Lo5DyL6jxjDsnIib2xQdwOPMAhHHS1VeABC0mKrfls5/XwqK9yH9INhee8
9P/Uj9jAkZXKdBB/ukvCDb3Woz5QpbbY8PochOWSDUeMtODgUoe3HfVxAO9RrobE
i9KNT2qh/O0PV0Zo7qSJvIHUc38RyXyJ9O7i44KU7SWdp5Xk55ZKvvI1wpK2QGc2
K4+vfSCNT6uaqOvur6plJCMHqvrtoyWnQRYi8a55IZxphtMazui3WE4uBHIKUrDS
jeZ8Dn1jbUrj++w/6vkYjoiF99CGaxPF8ekCBPCwhL9OdKEb64YyJVsgs+Do7YzL
xPHD5HKc8LTOptW3KtHHdEcTCjt660yEJ06iQAGr96sZ+lbPfSHdOB5Y/rW7r71s
zeu2FHvh+IGx+HRbPh7GFFf743qBtudZmb5/ETthHV9b4KXZ/eJVAW4jENgHklD9
YiO/ATGj2M9T43ay1zEQ/as0Yc/cJWBUZXwudzrZgtcpdHzfjPk9zChKWPCzVlVL
2YIa6cTWy/ikqbxY+KzBRUeKpeckH4Qluy84496qCg9bNvkRqjx1zmsPj/zDMr+l
82pWBUq0PowcUeoxLmVj+hpOHgtXY+byiMk2YKAplZFKofQV69sF2OkYyl/Si0hI
pPbMLTU2qr+i9FJA0rwiuVfSd6+FDJ9oDl93sS+2zVYATk1E6YlpySHZxXRrwz+4
yceybTW/xFhV8JFP9liuwbaNwJbXbVM/fuPUit1VW+0s0K4iB8lidqk66Sx3i8mc
xhyAh0N00+Y+xnE6CEcWZaTTA7tDsbeCvgXcx7n3agS1YD5GktzYrGONBz7+mpPM
lggk9c6wtBoKdkh8wl14GuN7wFL3QFcQVrvJKGTuwZy45/kpZjG0b067Mz5BKX2W
5+6rXtPj/ClXwvwnS0wag0u+Y44J/aPT6DlkO7yEDDZ8ITgSYw00D5OvOhB72nqi
o1G3AVvBjX7pxo40BKM6wwwvBVpG2N4NMXttt3JiOgdlODe1ps14VVZwH12NxpYM
yvZc+gCHiQJFpKwiDijJlZdPG9ALGXU7wkB2yLgNUe1AcmcvqqfA7Ae6OrhB9vLq
DDuuxDeJ6iHLB80aimspW6S4qfBTN1eJa3JVtzRdZCrFbsXWpjkOVex7VDtB4EUk
QEGumvO+t2pSEIlaTVL2WiiN91Pr66TodyHlbXJ4ArpJ2QrvtyQvTGTyyHhbMXBW
0Rs0eXDVG2QldcHaelKMqEKartMcuh53DknUx6pCFoBcXQEECBj92i63xyBLxteB
nwEtFM5GZ5Zl2o/XVPXB549CM3xRwxUiaKPQJg4qZvScEAf6TWfN60KddOEUIw6Q
eMi3keqI7i9S3aUdinQDE9Vs9V/w+SIHdUfCgwlU/VPWNJZv5gdjZK4oDtIkUDLa
5npj5ed5RkMShjFE0Ap2883FagqyW3qjWkhS8BzwI1mG3QJ1WHV+LnW2dDRTDGlP
fE0j7ToRTRC9yoGAWeGIwJc1I1kXO9VWHgECfWUIE2rFfYBRnljpm2goLaqXenKT
opglY/Z67sg0gVZjdjpVsZ3i4zDq8BwCn7qEUuccsOeNseAupBP7voUoE3zta1rU
koLHraHBHIlcfjFY7kzIT81ifLQlIr42O/HTg5zc53lwEkyBS59eozhzsYl+xrsZ
/QnGz6z48ml6bm38/MzvOkV8eyYfsgIjDLuNiRX0yF1HebRj07tCWBTD2OSM72hk
Ick7w4WhynNCbTp2DQS5aAoUGtKZz2CfjZEGd3W7tiAaemSeZSAfilVZMVqf1Xsw
ubnDHb1uk0a8I42+eHx8CBtdh8Dn7dRvu0vPUNZqXC4h+b8jN8jcp4+aAO+OOhgf
qkFP8ZRgTLL+avAYBa/Ettd9fvltiefV2d2+EFJ9m0BHZq/GnyY2jQlJxGc26ydh
QD8UlFrqXLrQBjfwREWQqSpmMAHJdiR1V0RcFRpoPRulb8JAsFNNnbJgEuGx2bS+
lJnyESv26PQ2Lqyd95hebCkIUL+JR7Hhc4akcel8/j3BeSgzmfKAtQA3Bdsb8LMv
RTzN7+z/35HRbXsrgF3w37b/DklW/5jDL0VoG82FHiIzgjEANO7ugaIVAoExA/n6
c0qPWj+CaoRIIl0+QIOFcNxpaLjxG3txRSm2Ata8DQSRwAsm7W5eMATLiYHm2tAj
l4hqdl5DVlyNc/gwz/d0LvfUp7ttOAeCJv1601a/phsJQvh+Aa+mmSI5u3q5icLc
OQAMm3QOhVVEgTmvDKRtXlM7y8nAODskEpBs4dVW34uj9b5h4j0jpnF/H2+u5G3o
vugE2jl/wrUYCXtHCHVwSb8Em6KbmWm9gzCjsw8+aglDoMaeYFvzhp/0mn+RoRQU
cf7mvET/EkkvdgjztBzZzb6kOwJfyic2e2D5Nzuob4LgN61az5Y1hzstwwP5NVgt
EmeLVDfpvtHYOwJq2R8c4ti8hcxPR3IC88qionhPFTHOerEWBk9NvPDkvNoo6M28
3j0EYjQFqHr9sMon8x8q6y9SccaHkqE6nzMcZyTKdqD/tMZ1VlMk80cZoawbKxy6
1X2SAd2yRUGXrWZIOITjhMGL80MFKOLkK7DBrbvF0uixq2ULuCzEykDtqpQrVIK6
XEQxU2Cl6lpyVhhQQfq7D+F16m5UpFciTxGWzBGbR6vt4kxdnPXwHQRkrTlLxEu3
rgP5xKdYmW9NK59tYdMCwIYfu/4IutVknMGBqqPYuUudziXw10/DPGn0TR9zEPpD
JdjyGdNTfBAn8Xe3W+g9ocd+mrvsky0XuSP70JITXxgl4UuXBTTTGJ9MpoD7s/7o
H0kkkuj9pkBcYcdPbuRyKtw0jRpRz9oRMoNyrpPezlxO4wvdOdlsNSlbKFBIF2Bg
qFqpUZBK/r+OQ1sQIKiyKftQ1NyFCae6eUE9a/Iu4Liz4DEl+kO3PLK3wRk/wX+g
aSRR8lKIfnbbU5iO3ixKzR7OczhqQizgkpgr83yl/EJGDkLxfrsZdCSnklAlipm6
AAO4NQq9x15kg7jUHDG9QSagWgFdF2CffH8tMPO/Hug018YqJDOxz+mfj/mKAV8c
6V0q3m3LggPNFt3Xsmk2Dm0TK0wdKfEUriG3ocHBxKcXGZPklvskeJH86ruSUwrk
CYmFIu8N2+3WTKtbsrVv5iJwam15VvQc7nO6y8Sz19U=
`pragma protect end_protected
