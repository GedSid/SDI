// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:39 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
plqR8+CG8tR6cC/TuraWMip4UR0O4ewygngH1rcuqfEsDBLuSbVjLiLhNQIDg36q
osN/K+BIsn6cPlxrw49NRVrZp1O6ENfRlOF2hgeBMOgABo9Eab6asM14nPeJLW8l
RX2h87AVQQmWg4wt0sEo0KFzGTs0F+qsnaq5/or4ZG4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18368)
XiY45h58NiGPA7KnHIBE2r/OuHfo8M5YaPZ28pF/Q6WXbX6PAP9HbmS07IbBkJMJ
2EhFmfHEDYJR3VcVeJZetuVP1hmB/pE0TLpHi4mpd79mD9YGrwdI5r+0f5SVOBzE
Ddp6atdUkTagG+lOQvpOkugZl7+6zyTh6VPTTwJDMiFd1ZtABraiebyyuHjFH7QQ
rNPDM2tKP70Dmz39R4wV3wgKC7a7BZfOyEXeCx+kvD2fD6tgChs/aXaoeN4XF89T
YhZjD86J0tf7q/b7eoyhyi728N4NmXRkQsqCHkoRdmtCMIoYI74yNPTzGMW69SGK
ylFIQq3JYxtgpM8Es4moZh++GbMMHJ9XCk98ZUmassv3LG5M1BTrWv+XY3dWyZar
WZIme7MTePZ7MXjVDgH2F/uq4tpZbEqyE09xMVB2bjKlXhZ1Rysc8PZDNTMDAooV
wcq4yI7nJcrOsEhRktsij49Q1bEfExSzthzkZEkXXrLvfRL2vw4ARBEHZ296BjIB
YNW7M0qYwnOYhjHYTPa4x5UHpUYpV6H0P2dbBFN93worde62aJePxVRmBsPi6Z/c
fqm3j5maDJBVddgMr3KLeUrZTH8VvG0DARDDvvnw7MkK5iuqxndbUy9ieYs+iR2S
WpIb4+X2bSQfWN/ajhQGrTyRSwpiYNL3KBSKkS0qlKyRGGlh0SDwEyjK5X4R2Ytv
NAp7TC55a5CmVUinfNAKF9ATpI+sC7aeur6q+iHjy5a7S5XZfxTtS5z85nKnQXQg
nMVMEe+WlR8/vckX8bPTtKQtOPRB3tJEl76NqOfI1sb97oUtZUoHaIVOOvfEKSIt
dhA3aNOS0RnCMFkgaihETA0v+sXh0t0YnnuQAS2jx0dRPc5VrN07Kr6L+yU5Llsu
hKebCrby09MqxUsFG786mE/sA08gvniYM4bM5eDDvLhd+cRo1c2V7K8hEcpeV5D0
QaJwXQ+2ba9IAot8Zv3bkGJmbkiWgqZjCHDEDwOiz5kDhQtYrMDDAipFl+K3IxPY
G37ULd9WenmgJJlQbe+DxfvJjdOJWtxtMD+tV08+QY3M0d0N4dD6ctIzE2LnkSHk
MQjrX+Ra0AYc49JsucHQKvcgSv4qCWAmmlNG/hn/LRsqnsjHobweSFZsn1VAb8UJ
TIBW6ulUkk6wwNA6yGa9Wnd7WxEcuJ4N9G9ZkTACZLVCCCaqoZY73edXetLjkN5M
bZNNXYFUdcmhBd+EydIysSM+VeFUCDEUuH6OIT1oGXgYmLJqCVMXvC1yq+Muvsop
h3zomsTJOOnIsPpF3VnWExC8NRxmw7kso/313Qwcp3kuhJOY5vJDLJ1VdVXCnAaZ
ZJdsN4Hax+8ia7al7o60bewDvxtywPeZ9hwMSmkZUpeJRYpILc0Im/bzwxFizIMN
3kSag3HoSfd6SEuR2X+2fmJHbPzhrVom3mDpeBAlzrivlxnDqt6btyOizIBSQ2h1
6XOZBsvGhFo344qkxiYeNQbjkARD+X2XYBwOY7QdOXMYCmFKWCtgafWjsUX/MS++
HjfMIHzBDNcS10FB+qtYPD7u338ynzTEEGoHHqposCDzLX1y1ux+i5IYO3uJReXx
Gqd2ZxEYo0gm6a85/jvqN/IA1Mt11IHuuhSBX44bL8wRycdirD1r9VHs0iUHWD3b
OPQanCNG9UOEUHSzoJL//+HxvGkTzTKeEbL5Ni1xcow/eZWpsfQL/7FbqvuB4zvh
7Ly2sBoJd5riMhy+3wvLSPd3i4w/8eiKWpU4wQmB0TahGGCPlyxjfpBvM1q9qCkL
ocfFs2uuZrNQ+hU8VZ8wx+OnP/mc1PN3JQCjtU58AUD88dE1k4Pybezwo8q7C2jl
WpJEhRwtqOn3pg8xc4LUyN0G3iTOLGQBEzLKJlRQn2gz0FQLjFUMkmh8C/xgyvcb
aSdonNdojj3Psjy1HsV9BsUl79izjOGzRoYNk7KucBrkZApvGo6vw67/QPjCJdL9
1il0cBwhAYFqjPEwppJNGG/n2v6oun7qSymZ/FqtKDQQLK3GtXoV7Ep2kTaqzDNX
Go+dD6cH13C9yco5uR4pki1oItykLFlRMbHSffwVUs3hl/Hl2SI3CdfXW1bgOuqB
+9iAEH+H0TdibIIGJOu2AyPJGT3nOXqq0EC017qqyrZg+D2/XsbfvWhydATnwZ4t
TJJJHl9tTc5Qo5sGcAKUW0VUF4zf4P+XLw7rN6azDAL5h3qpTLyvPUDxAw1PSHtJ
Dc3QNZAmTxIjAJZoTH0h+lygOiziEjQwDLFZ9n9FSNu+eO16vzWF+NZXE6IW7nIN
9xLRj1tu7/Yz3hUT+UFasPqH4Wix0oQNW9qlwUfoTLHo3QiWRqLHczgK5CP8hWiF
sA0C89snqzxFiqwvN++6qcaaBuN3EtpO9BxutGekEFGPjcmx4uOOSOD0Z+W1sPLd
6BCAuVXhggCrHN6kFpFNouuOBnDrbFp7UsKyhf8EgedbhT8CBlUq/WErI04sAyFl
6tUnUdc32HStXJInMTMapOmofyAUS6CzquSv2tQN8YmfUW/HfuouEtQKdnu2a32D
e/bxs3fbko4lVcxuith180snoE/y36dygQOYvwDCdego8bC3xYmzw8X51AP1FhQ2
QyGECQljk7xmVdanS5lz3dwE3qHCIloOzwQsHyqTjxQw6c9o0t6oU0EIg4cl+ayv
VYgYZNTAFgy0N0vZ+x4mLwocUW1rP1R9p0Xff3K8flofIqPmqex1d3nPyKt6gzWJ
9XPTorGsGnjRy53oJEMPpwOGUdZi1qi+USc13hK9HWCnh9PWZvzBRMERBwaibcWI
Nbv18ncHzTToSGXtzs/POdvjySu+IVFZmZUixi6nW6S+K1FDKgmXAmGJ7k5vY4PB
IFHWuQsNTuPBY6gaDmGt4GmNilvCXF8KMNuAWXjzV5RIzOamPSK017EXjxPduI32
ZA+eGhaY9EyyuikIiOX+JDCc27S1OpBaEfjdYnaLRVuyfyXw7hTWX+sXb5JmkjaT
bk05XI2LMHXVbJ+VRQhXu57I8/s53K0dtNXnVdkQ8TdrtLAHWjKDZ3ZdzUsjtntA
GNpQMHb9M8Le17cmM8wSuH8iKwsY9mlFCS8LhQ2IIz1SAtPJBx+4ppC0LNAkYYpf
AOf1crSbj3cn6zua5pdmRJSPiASfl8zfOG5h64PUK68gRciLQaOt1zPgqaEd2vX7
3e/HbelGQZ80s256r+/3hyW1OqXbyMoGGzkDjWP/WdGMXx74lHVlncRcbKuH1Bdk
4wLlhA/fmX7qppN0Civ7E0JHDLniz2fRa4nXkEn9ZdRtOrD3YHohKVH1DERj36/v
g1C8GFquZ26Z0u2prldDweRQvpMaapfaW3WSOroKejgfcqg0gUu1i6wePfSvUhtI
GqNvptOE/N5R+hbcPYIGJekcVNgTcv4gi56IQmPoj3K+++3HlsM1Dwopk0qgGUE1
HFX8fudtfZmqf8rr8tWwHDXiGUGMggqMFJidjEB8gvarhUkEDs2JML7uUHD4qCTq
Kx0zVQW1WKLk5UiWHfBSt3mLMmCqtFjv67MqL5mlkWI+RqQFXb881x0GF7txyyhW
9esRNkgTQOV/Es2WkUTJnYv2w6lE3EBJ7Inmut8bxBCmT7CzNlUu5UdE4xmuAYIe
ZNXBGg+ubzD8/Xi57CDK1n32sC7tsknmfgrGVjkUeVWBU9ILtMhVyCZq4G7GJlgw
4fPADeZ9RS+kIHIkDa0WH95GiffZd60xKJSotUuNU/W6IcnCdv8OPLnAUUqaGEi0
zArFYQ5ZEO1I7kuy0ocnNGAxEDM9dM3pE6MNwZ1eLyte6hIf8P/x9ES/XIeD5RZy
dBSmr3ZniIbkupv0Ujdacsee94N8d07ubyRWbwhOLHYf4z6BSvzt4h2BrwlZKZZZ
AKmLgMM3n/VFClyb2RwklMbv7piUcRgydKqIE8pmY0L4kfEwiQ4heSSUN/fViZ+1
hJs8STNakeV/kXCIVdZEOJchDI5wd5tGgKNEUaEsOivS0a/h0fvJN+NaGzB0M0zr
h4uLkydwKAY+x+SCStg4CrUhONa/EPLt+5658/3hz1tjkcBWKKdGNicZgLdBAanM
+C41AM+mpBO6JWgJPE7nRdJx/+eAFEqPaYds0lowGzUPDeraz8J5tP5OrOvcMx31
sFwaweSik+55mVnjjrchSq9HisM+Cq/dNTtWgU3pCZBSwrZ+DqBUT3OLfVYmFj+t
I32xJOGlb/JAsk7ZpXBHxojNLY0vjUXmpimrjjXQzwaPRBkbzT0i+Ot59wpBNXNs
5OjpEIT9L+KKnTrTbSFvNKTKKocDXuMf891eYJBImOX8ZPN9xwBIPyVMgETYH+sX
8tcd4HhRKgFSvwlYO89Jxzaj+4NNzMipry6AHcI9Mq/izGjZsJEY49WvW6HMHQ2e
GMeptTkesPEtRZlzyrbn82qlahNqTVKwJqBLDRT9F7KzOaHtxHxF8EXcQ9hTXmYg
7xNylcZloMPPbIi8amEPdrV0Og5LtZjeF5TKrH55vRO58Ht6jJK6biGCSoThBWNe
ePrvYR3YHjRHHZs890b2DukuC+MU6ZzqFjC3vj+twWM7VEsyscHCQBlu0sTtopff
MLkXD5GA6O7hwAzu23e1HD2BjK9FUxPIEV/d7jsPZ3lT7JJ2R7DfVQB4OjMzBP42
vGYp4lsqBd8o4kRxnebpTGZ//o69Zj/ocOWlEjMjtnsa/Avrxemie8WlvS3Qbsre
bTNEaKtm8bts22nRR7krDNjDokGNmnp6fyTYKzwHy0aWHffjZuCJD0A8b31EeRC5
b4raCp9pv/kF9WNWlvhmeQB7lbcQem3+J9SZQUdgDvUaeE79VssoYhb6xNSAxWuF
orfgdV+ICqkuG1/wAPJAkW951alDOcuDEctQBUnJS3tNOp/ejCKV0IHvEDIFh+Ef
iglY4g7bYDxMDyZu3Zbt8CCzUwAWPdbp9v7u+m+O9zBDptmU6SEFcXuZYxBxIdfd
IvsgBjq06IlVOIvXa22nzt5NXc35VDQuYOdMj59lMCQ2Z5UubKgaDkbTkEE6Zmax
YVFdUNDPPJljCoSgncqgo5YAEdZktBda/56QpwkuSrllInirKhETRsG+MSySWT4t
ATNAEyMrvuHwB0jCCqh0VmkuzZKpsTxw7/TtwppyBW2D/ULyD5PdBQJForEfzB2B
kpMnw2dSOBOsi73XB12F0lr7NtbvVJnV3nxhvLkRky+3zYY9vufAuLNfG1kNeo7M
09jWSEScBlU800zSrDZKuMo1fkJjM4bT2qyZw5vmrG2G8b6YNVxoWbWEUcVTEnWf
TeH2dTDAogzxQTzoyf3+EJg3D8KItBZDN5PbYwKVc3RBzkC3DKDq86FYwpouujZx
oeRyYHEZb/47fHJ7X0mSwZs15Ji3WamEmbyN4tovSz8wdpZFQVnLtKi945Ed4qEI
nX43os0jYz9Zpm9k9MPMt3TWPys4cgCztXw8v3/qvycAibnX7C+pwhec54K8zzIV
2DclKkqfbR6llo/FwEWYl89wQ46ammmxw2A+Epw9htuI+uykfFxob7CyPjjdPcEN
2u/i1QGpudeCWKkNoh9Ohska4wUfX3WGkYf7gN3cd3dLG8tHZ7k3oEZmLIgYD0F5
p0MJT9w6bdUIlal5rVad8Vnf1ASXbaArWZGQcDBrbikfvYnVsgVA5ZCvcqM12mpX
hVB0hEi9zpD0Wm/AOIugp3lQmB8rNBrzBg8uK6arkvufT25BDrdc2b/3QRXdnUe7
RqLziKQ0SuF9RsIfmsH/UL9E13bKwJOaZJ/DO2fv13rPCIMFCq6c3TPszuKuebRF
5m6CCCeFxRufQSXR361/hSVUHFzrsQnMhUL1Mazk1Z0xjV94XxAQ4JvSel36RMw4
mbcqEL1AIQQIArmbkZS1/2WQrQ5kyl573nQpS/bphpp/Hn0QijHCt0PhdTHiWO4W
joWlWF6EI2KcqZujmH1FafDnvNhiisny6B/xnS0iH3XrJWyznCMHja/3+qiXoSMu
ycHrdAVSAUzxT1PyUjmj6bfjaxlyGOmF7QexxjJmmR0r4C3pk8NZiaKujJ07N90D
M37tMviM4q04f7bh8U/kod5hAkPRFKqb0yVsy8VbPCRYL+enG5G/DJqxW2LZsEys
8Aq+D8RWkZipnHFB5gNIXAWLgKo5fgaTYVd/qQTKA6r/FacdmxxnhgZFDUTk92aO
xeRd83HJpbX1voEtXxMcZdkvskAknsdc69fk31bga5bTzXEnTRMMOrGREXDfYkrL
ttxAJM7OiD6JQIXMOEmbUBUQ2FQYcutV8NtrP6rbicQyN2Mmc99SElw6y3G2cPQk
MIqBZFdERI+ltV5GQ0W4s37pJj2YyDOIG+Wa3P10QTZoPN+zQj1BnR8I+vS2cCj1
Ru/GSgVEY2hWwMvOLfZjazUm/PXp8aKCH8SRyRj46I7O7/eY9AQsUiZ4JM4ViIWM
oaVFMk9t/00aETNd95Rw46CNzhpvbAWgjVkGmo2lF8Cae6IvNZBh5FAPpo1Ex3sx
ua8k7jMVeqg1Rfderd7GNeN1b7F8VKqlQJPOKzIEpjPTXSnRav8N0Jjn7cYkQcmY
eK+MXIahtUnQL0EM76Pk4uWUC8LfHnW1yqNwPdOlcDqIz5XfU518GvimR/cgaUcz
4fCwpufFT9pcrIaVWdSLG136zcjdFAuvZZFU+Hct1V+U12igTNNuJN35PHc5JFsz
Q1ht3xpIpBwxhyyFJmYGmSHepSGUWURiZd4TaMUSjVattcCrd2QUv/4xIp9e12x3
KVcN0uKneRk93XX2Ei1Wti7vbro3dgKoCHhPsUAMn6UBF0Mwt3uVckn8umD2NoG3
Y3mCJkIhenMORnKdtOG3Kq4qm9bW1qMVqpw9AoDrK5Vj8yDSj88vfoZLMKZDiDpn
1maAtRKxLPTY5didjZaw5Rsb2ABlCbav+pRad0XuU2zwr6VJ5yrS6/dPI8jNJbiq
9CYBlF4GIveLIR3/iAaTIOs1vrFjs8VFcw+qpthFFNnV8NUE99Ji6as8NklvfGr/
+9siA6JfwVPCocveFuGAFWOalfeQKXOTuCi+iAHqmDU8+7h9VCUfY7MzHCRPH7U+
yJPCGuYgPXC+8Mpb01W/7ywRpaDt79eva9pLjjBIIllunc3PXrpz+NbSdtkKGAiq
R6G3smF4bYgGIja3ZhFt76ZidlF9UWT8GOoLh0bxe3zXPFuoE7M649WR1x8LHKTT
aUoz74f/87TXENmnxeTiuJgug+E5fSH8rne/xABZejbrPwiJmxPCCtKruaEQn+83
iypj6m2GALq0WGXccICh+/GluF229wNxQoLOO7d/Q+wBbhzPQXS4DDICf6GcafTd
4oX5vF6EGS3b6pmdCI4/WguykUORoPLF3YKxn0c1epzgnMVQQBiX32lD0EXfEgTp
sRMFpOEScZ99SzNWwpVNK/scYAXuoWxtsE6g5GR0L8ILK1oL85VqV4BKY62yJ51Q
nmrQMR3UbDVzV1eu93ad4dZNOisEYBJ/KGNNgixIVQu2lUQwWnvQkt3ddCPqhopc
Pc+rOzKhs7aot7jDJZDbj2LT4MvF0nU/6UgR1o7P+1RRluB+BgVEEwWWLf0U1HmP
vy3m7WUeSmJmZZt7rjneiMgHIdcAdD2xA6OpurYW3uwDm3/xhJ/bnymD/kRinKPk
pAp9s+ilUEXAP6hVNHfsuLQNFokw1+RE7qOcm1xPOaXm5xetqzsvAzES79WI/ARu
B3vdzp5E9GYl8E1Bba+8egGEk9SGQaMEKG0XLllmQCqL1u5G59wUt6iAQ0Krqa9F
h9sbzwUs0Zy2nDzIKfyxMFXhfs0dCXx4F0jvwel2BUZeIv4+MDnuX1Xhdwph4Z9g
zeOs6cU/4h88ZASQa9Mlq+VbbI/tNJCN2lEAG2V5gRftQjDBjx0YYPYCcX8Ubrl2
rGerw/xwYuN0y1XnN84j4UgGHcvWzF4C9rhfStrvcfv/TfpnmaiTYWh5+/8IJCUi
LqsTXfAZW4RdnzEae5guV9rerTpS9jK29CFY/YNAKBGb+5NNLSk5YOr6SNzdSNl9
+waeMoMJ2BWrRUZs5TmYj4vzY43YuqlZ27NIJ9ybnZpU7vUB9gDO270IP5d+2ksR
vzZBfPpDxGrvlby7J76uZa5tX7wkYvqC1F+rNdRaqb5PKuWBeBbOp2XZII/4IycD
7der3OF/kJBQ8JjPAurClOrRaqXwVh5mvWzU4WR5VBWP0U9GS1P3yip8rpn36noJ
Qr3tCZld3m/mUMMjTdBC1bMjTIVswGq/l6yehB9oUwtLZXpR6dUwHOgNj9TYcAbf
vi/nEqs8LDDkTvA4mK+dZRYDWRwYRnF4XRGBY1sCbnrFS737lLZ+80mubMqXbyvF
U62Duth9lAXp44Zvf3kIf7OJTR1SjhL9IEaZC0+C/OG0Rg/hiGbIJs5eaAH+xAuL
F9Vtm7GwYWxIEZ79jKjM6ymMpBWcQYev9f+OWWbeFDY2VE0cIm15raAa0Bo6cP+8
zUj+buSAZrdDmbCduyWr411MqKrr8kmbWwVxkKZqg3nYdo5U72At4lHcJ3Qk2dwh
afu4fE2rqehvLBhPrwMeA/b94sRH0KzysRipRKMXxFMdDydcnQUi2iBVPSoyK5X/
6e5VUe3hK4obkhpOl3+JYvwHHfFL4D8tiJMQIcaysn0uir2ci/MLRJll/kl9X/0o
3duqxcapspRpnb2faDFIUOrUUsNcb46Rj3kF9YcSgXZ5LcXryaYUWoryD5ep/4wk
u6FAebgMGGhtEw6lwZTGjv4h3NabH00XhTnSfou5HRBZHSIxmtHG95grAyCOcvUT
M1cM+/lnEOHVd0qsv7Hp0WxZtZysz1+7CHDydKPXkmRcnzx0CTaN9ZzEFLk9mrvT
T//r7zNv3DU/mPBwm+5Ju4vvZcR4zOvwcmOV9CTfwLxNp+To/0Os459p/XbulBx+
qEIRbgiDpOQDVwbq04CHz77tshTs5m31cgoVrQbC1R5CwVGTu21KQ+YYX0FZWwNX
94ClYpRDV5ZUdFharK/zWRiu9yJy8M4/sLHJG7kaVlKmcokF2gO1/AMo5J7sY7Ey
u1zFyPx1qj79g9ZNywdy/KwO8PfhxiLBAyQTgDkBU4xFkg4NOQel/QJ/Zj0Dkad4
vrJEMA5NKDN5IvHqYLYdFBD4tYuhyqdnryOQ6U/KfW0yX3uxkNNFoJCUZGn+p21G
5PCPNSKG/61KOwSRdvJZ4nSwatlbyzTQye+naOhlQuIJl7HXRBsRZ4Ddg5s1yszn
tlBnFqC1VJWYUzOU+gFGhzjHziBmA5ZsxKnVVlM21ZJo8HbfF0FiZO9BQhnv0sO6
+b3iHX/x0vR6/fWZQ0kiC4KtKk7ZScYmUjOlhwcsThb3lwBP+jchuNavNjIIrNQl
StcERjLap9vIIsu+MBv7SrTi8uXI1qJT39amcaN4I01axKafOzqaFvV5oK3MP7w9
/Gf8932d9+HNIFGCBAOLAJN46JUmIv4ftTUXbyLsdbORByx6vD5xJXUMjLrTm13l
umECTUcV/HWtKCg1xkIJ9tVkVZFSHiY+7AIMeZ3wb74UKSE2gsfbp/hwf4MPBh0A
A5nFT1wXTH0VTZxEYGnmvy6qrL3+54byp2sTB21WFYn+mQF9W1FxEF7NSuiDuOX2
16btRyUpE7evlswUdmf1HUxp+ls9v7arjk6BIrZjrfuwuyKbTYapEh0HBR3JPvcb
Lgz5Ovs6ZqWUBvEpDRNxVhC197kqTeL7VpKxxTAZBSsU+F/c8IKWVmmW5KbkY9/G
UaQi2n1FLAD1MyCcgPE1xRNmaGzGN3nQDu8BgYvmJvRGrAva2x0eJOQfgCQOMzZe
Lf37qXd/0zgeYMy7fS/KOBOJaNQ7aTo0IFua4MyOxR4pGZ6z0RxR4jct4DxiDIkj
64Le8uBs6wBMY4L2TT7cbX1rkAT+cCkOezOBXZKTUaOqrlqTyOJ6Rp2tH8/gF318
MKH8SSnH9REPOrY+FF6W2LfDGToDoEvBucJa9mF3hGKE34HC3Uji/1/i0FJOKa9Z
Jqi8KDmilv27vBt3FM0sesFNKVEnhE8Jo/0OjVV0nPVN8h28kojEGtR1rTZ4LrD9
P+FhPbZ9Y8NU1oEWWN9yaAqjShEM/uulXdivb4ajqgUhdJD4+vSZT+1IfLer3brH
hdlMJERhnhEB5HPKBD77pA3wZQjZTq/bwz7HG48hHAi3Wp0tJHCu2i905dIgt2Uu
Hx0sfY/08KbmiVS6fPKT2Xfn6jD4ZpNhSxh2Tw6oCO/rXC/1nOmD1UpAgHysvoBc
JvWv6KhMcF/k8EK749zV1D7Uvsy0VSKhwEmvshxnOLLaCBiO6o+G0XmHqS3UB4M4
RZAskuEzqtzzDaw7LiDMz0EobfoYPQoawEjaSX4Wl6/lIRn/qfdJM9Wa90YoizUC
zvdUjRnn/8sLIRWMgXkWjGMUmkvq1iS2c+BK6VXjj3XL7ecrVbEP+DWCdrTbgI45
GmYG7d6pRsvvx/9gO2WrY3PYmhXHpoHU8xtDUy1hWj0PiAOVlyPWWrW+yiqBRnjN
RQn3NHMy073D5kCLcix4ktp9XzpiPDBw7j0+LS2bYOzpXH2nMZTFYqKpC/OdoDVd
g1+F1kL94gD7V/Af/URyosFaubq/XaDSUqk6w8EYC2V2gZlNYuh1c5m9p75rzumV
sdxogDikQ2wQROXk/CLx0u4cipzH1txxvHbS4a6jiILzSXJVn5Ep7jJ7tZz/SI3K
cl/3bJxIB+Ej5Ai+S8zFVOcBSgGy4vgY3rrEHDlIlfPXRmntKJlFUq9ZibgUEnTy
EEj1kbhqeER9hABP4KiHc5ij0F35clVaNM39pq8o6MAZ/Yel+ZTCYMdMLm2sNTqD
aVi9M/iW/y3OwpfajcplcUVzuJqfC8WkaaA4/ujg6wq/Zh5uyGzVvGe+mo3ZipuH
HCxOtOH3i2C0Egkik+kTPpmmc8PFy7Nl7UFJ6Gxxq+BnYmlKIuQILA6CS3bUBpKr
f845ImTwvYvENHy0DXN3Nza7K/Xa0PIREszRhadhP2++NmdBfuKg46M5nr9Afh7Q
zD+P9US+XOmvkHSceJX151uVPQ/N3ysNPzjlDNhkG8D77S6eY7kkYvAfqvSvHICi
M1zmPX8EBayPO32I86X9Ehm7PY/qLZ8R9v38voeWqJQInVJe6tebGEAWl2WjE78V
7x7ReulT6ULW3ICcoPXYtWvEsmw4kVwUvX+XB7McnP0qgv7WIdBV5pB+WtRxYh0M
YuUCayWOpvfda4Zelxq3SS6uIVdrTraTWsxZcbWimMYpY4kL4w92NvW+kr75c1+I
27FeJIiQjcQUL4CvBUFHiIOCnSRG8UTEys5Eygvprk2+UGsZ8TgSE4+kTCzl6u3a
XsbMhB8nR3fsif1O5JpI7BwxdOwWwXuYdkp0uyTo4dLfcaQfjThtRWqgfTLD+UGL
mA2xjPzBC7MgbfW703R72Xj7LAjP7E7uOV+N6H7fdx35VILIQvVJ0nf192Cz93GY
vsu6185V1OmFPFT1v7K1RP5ndKwBxxq9QzUtQI9Z280KkTOqtUAnHgebIY0dqq9e
L7f+LuCNkv3izT8s90M25lh6UXfJB5OCzhrwbD9BOqI+CRauqZMtG7Jmfd9LLhV2
LWEulHolGGRvLgApvZlNCt6wMBN3gKJrml8mVZAYeHnWAw7vEJZBSH0Ynq3Ah1TE
ksT0R5ZOeUfqg7ijJm3bKfZNdaZKiNgEsK0nGhu3eoF0zc3BSbSzo8a68Mz6yFfK
uP5KpzRCt/ZGRZJ2WPkG3E7S/yPuTPWXjr0AbWsQNILNTOKQArqOuPlwWBVOhwmX
vbh/pmqz/BKZMEvUxwo54fOYQ91lW3wFkbn/0Emk5vC6gYMBJGJ9a66GulnxBjD1
yKjJO1LHvi5hDwxpWPQTFNa/5JAlySjZPPKpuuX+8WUUKcF/haprpDmJUut54YCm
Gpmz3uN+WAJxxokaptlAtBZR8iPgIL/IMp+6aEktBZqd0syGzxVw+36yL/TZ+d48
HUdVnC9hqG/kC6JoCdv3k6pYWz/nB+Jkm+rdJEqvg7k50gA59Sqs+5ljfoUWqm2G
ttAu6h/n7U9P0YSJ2hUJrKAMq4ijhO182pKlDL3pLkJEZ8wRePHIaKkb3Eerp4YL
+ZJFwqpvNQSa6mL6BPfX36Ns1hGt5/W1PiXsLcDTMSdtn6PpLM6gFpEozb3CS/uM
p5ovF7vOmIRexPPiUgI4ct33YUAvj1S0Wwkff/SzxGCS5V2y8AmMnXCRaQpKqbkz
UqcKCKHa5Z2pypO8lPnVAoenTfxN34JNQTOxbLi1igD7F0s/6u4RQ6beuHSOCZ/B
2dhs0KSDwR1l244q9KEdiat4xruKXkq5CNL1Cj75kzbVJO5YiLEPn0UJ87v1M0Kw
cDEy1fxCORx0d0mi98DmJaFBGhBaTV7cw3JmqiqoRVgMM3CFO5p8a3vDcho12nSr
wwmgUkOhsNxL/EKQBFK+hT6EHsUlGJXumCdZJwn/O20cQJareOiMoEOO0p9DzYhq
gkfX//IR6eBw4vSrcEQc2pTLmMPHVmujkjoChDKhJr+/vX1d8coftbDLiLq7m1nx
sZvP1OpHOyf10MznNu4Hbnii0Tdmz2ZB3xi8jgvkF/kEWccdSG8/xHrdnBrxROYl
EebzCUiCcWiwOlwpRBRJcKTnCIW4s0R/Mfi52eFtVEkV+u3F2WpoG9oM7G5eadA7
pXlCla1CyBoOfrZj4hlyX6yl7GHveRe6c6UiLM9/y6XjueX5sPDjbR/nqtDJEwfc
1tnKX3hkKN9Vaz0jEjdVh8xHRx5Zh7i1lw3crqdwa+eZFh1h3MgEzwGziZs96NxD
1EfjGJSLRZq66EWEAapXx+sn576Sidt9rTuXVFwBueozp0i3ZqSFSjGKG/ZbQlsi
GqjeoUPNibsZYLdg87qRa0hsL6H58JDp9ivxvVOGbCo98v5BqNSwRI62DcTEvgOS
9GFjLVMX5gyBC2OJgqIK/0+pprPINobbr/8+vwTDl8FBN5+hE3/RXCbfg2ZXr24A
gSnpghDUBikZeK88MCOMEXRPLr129I7zIY3SipHtppYWV3+kfNAiSdf0C950iBM8
ILSAYqsnx2yEqC7ldbkfYVSgNgwwga8uAK3PkKVHYQ6BA/8tdZKAyhq+xAq19PJX
5M5+uqAFMC7FayaWGw7CLHNGlau1Zf9u0OUJMxFPn9uRRWE701egW8bw0WgtfNtI
ecUH1yxlY08MXmLDrsimY+XxC7EPWsZTFpWbNmxCu2O+flayjzBOx/JkCyr8XDB+
r+LKlBGx1HnUpdQklqBvKWW3jARc7SGagg2wZLZ68dfXcs2TxQ99iRDBRw4AHXCj
T3jJaYgSxnAClK0E0hHma+SE1MMvTHD85eyBWe7dFEOQ1ONLnubEvVzT3zeq8lg6
u2EFxkkg01x4OXQK98vesUJuOnYaeYAbp+auLSFZxtQ+v5ZvFqyVWkJ+Jfr3wZJu
vcQAInBpqdefxzOWC332wqtcxv3BKVRb6u9OD92aUrzBTeGk/ZKnVJ69uzCzP6de
ZAFprJHdxw87XgFXbaYH9ctIyeK6ia/8BHy0tySQZ0/WEum+FCdLEYDyF5RkfPsF
0oaZ6d8XfT/kl34EQ+U3GemI1Oa36/1dtCrIPICQuv5CR1bsL1Q1vdNRsi9vkYZb
tFyIJqFEZIx3t3cU20p2gYMm2aPyFlRuk+R1ZYuqGoaFw0WDXU2UDvcvomqemegh
+h6Afrjrnb+XHSzV2UOrhY1xx9g7lDC0Z5yeQs0bNjIODNl+PAVWsPsodlWkUV2z
PCppnSr35QypoBHMQxXkYQV88rGXPMIllJWXMzSDPL/A+rGwuTZb4/DJ7DCeA3+f
0xa7RKC6ImP5TBBgUirmv9HDjQaagPANO3W7d+TO4CFB0DDUQERKyVDpMyj4HJU7
ciXHFt1p5vUIsoyRz3PKczDGce9Qx9GpbMh/nktTelwKnP98leeDf06QXU9T1Dv8
/FDHhvNaBB36QdzmgbOvW8yGbSfwrq07AR430kv4wYqh6mxQ7UnIic3IKmu7YdrD
/KPllWahwHVxi6Vx6vD6Oy1sPDQP764gxI/1LabFvsUsJODOO8ZIDl1/NIsZ/XoJ
grwWJE3ahWE1058H5dyaydi/ckL2W/PmoZ/0g/21pWLDPQGPlJeC8R3JpswZOfc4
75khx/EDTOwzI3ynKGz5mwM6JfOpadg1pShXvRr8JQBHQrG0BymN5hiuGPZNYY8K
3MIb8rUsj0wTXFv7JHNdIdb4jGvY2FoT8Y8JTPM7tJeD6hKrNbKeu5QD9WwAm/zU
YXhFaQniabeyTLvD0MbOC3rMkgR1eOkFk5lFMf4l1fd6v62B9HLnNMEPoKEJGT7o
LepjUriIx+YNlogsNxVpJS2rU3T12TpsMwgBHK7syteeGPMTnZYQtLHvEPcclGvd
OFWOEhum8qJoEFqHc5GrAi1uPylPEZGMvKtL87WVXdGN4zVrbKCQctrLgogaRKYw
pdKnstnIczAR0TmBKkog2TpVhIGhLo7G8rBsd2JL3OozkkKjSdOqgOrmWdEqT6of
3/HKlwmsWdfi17e8uavkc2DhIaUuQEhjXPTRJjTnF5b+K8rMZE8q1Hz/jQ6/y02K
+wowBIpox8HETA6kSpIK0wAj7+I7gqTsPj3nz9ipMXvHtX7yyaPvQRjtL78rHAc7
RMH+lRLC4Fg7u7J8yc0st4ae5uZdAUEmZAjKXfjdANnveVHvqY7BJSGUeqov5SM+
cKT1J/NBWYCT7ckH8O0t96MFUmYWBWQNm4d6ap8fYzolTJ83c4TpjQeKaxgzK/S/
wLCR33YxC40F+eo5bTdftlwkzkg8mHcNCQawUWWTmsUW1seagV+b+CbruA9RBN5a
hopDnDkJ0cZl1zOOxecX0nw7A2BeSkC4FprSO6wRhWtsQJxzYJIOw2ruhvZannAW
ljOx3KXYZgchFmXYikOUmy3yBRyoHr1nz39L7jOG5pHc4TseCOOlQdMkVJSbOMp5
rTMd84wn1YoxAHpB3DjRXQ8fm/ZBEoFFwOVodemxE0Ps56eDDryWeLLky0fLQy06
ECNnm3pxH9giKNYVvqCqE0ZcZBSrlqP+ZagIpQ/x/Mkx+sbgrba7xeaKzGnA+ypN
Nuffnd4E2HbVp9WF+T7ijs3c6RcF0fTRN7G8y+uOobFeUK2NCDHVDYy8NIkFElcK
Gq9ByCQqDrPX3c2KTA3Qw3SaRx56HSShlj9d2yg2iSmLOLy8YnFUqX30cVGak3W8
th9UwK9DOXr5C8M+9BBCRGw9MaFEziAf5aD+z2fg3/9CsH/tgZKRHltCGvobsEB8
rN+RbXwUPszzfBuYtfNSgTQHqg8MXzykTPJDPBeVpFHumYv6AGEKP8Bo/v0zonF9
a2eaeEdLanQrPqm+BZekulJY218tXEL/QcvTp2X2FsPZ95nrlnhdSvnIQBV08mcl
LakQKUEzZKTj1lBhvSzD05DRbCjntkNBvMMFJsC4opSbPvgMQI9aTCdpNU8LBkAg
f8SGwN6ipjx2/+tdTRps7egGUJfWF5FEzg0AmFDD4HEaqYF7MG+sfyKGE+m4xw/O
aQrPJ2yAmyfuCzj37re6321Vcb0XPvoYonmtYVtWqs+o95qYLsRhztwFJU0HJeUc
dHaYgBonTcfQTk2Ky/kcNNYNsyFLwsaw63m5T2eQnCx9SHnCNFDadXylWKjlqQdF
rV2GVc7PdnuIbv0Ff2U/jhAzt73Ao+V/UontvfMN3kPQqh3s+TLSCS8qCp+4JMQn
1YUgnmnO3+SpaYJnKOvIY35ZnVgV9eh5tozEo6H9zg3GjsWJrkb0kqEum8vrkLCw
WT8e/m5D/004R1MKSBIhwvgQ8MLBeuM2MtWpeGzqtYeGo1hx/pqrKiK5WiHaXcZk
FJNKMOJ8IjmmrexEtpIHBEV7mowOcLgGQWe1COaiBgSVLyqIuLhAiC9d5RmgYVod
I8fskzB9cFvHnEHSWpQgvHZzUlVt0PbZ8cnttZLcuTruCxCz/dOZLpX3Gy3YQM6T
VGLlz514F5LaE80Y9jo6FLJmxdk4OsCZvkCoQDbC+5FtpudCL4/rRpL/Wd2rgLq8
QKYBNMNXkdIQZshm82nYl3q9uM0fAOH0wSeQhfjOReyRE0YsJERhByrvdOS2cAHn
wxrl4uwvD+I6vdtkJxKBkZ/5gauG/CPltMoDtXXlHl2EjH4Uif5Wxi1yav/mGoIJ
g2CYnUR9Q/WH+IjcGX1CEzClJDPfFjNXnvJmk1twegPPJ1sK3cXgGzpS01V4BDLx
XJ3v53QcJhOlglWxs4rFBYoqAoedh4AldQXpfmQTS6wqMchM7uvccnprKzT1e8CM
hqyt/I8AgAyNSBF/MXE3nSt+NaCtfSGsmS8JFvHDkZuDXkE/iGvi5V1CF0Sgca6I
GUBiZKydE8FRPR4XMqaheMajVTnHtbpI17W3iOGVu2KVRwMa3Q8rjy0VQgnYSoMp
BAmUPOScCXm5VZoCBPa4tQFRP57Q4Cw8T/OSBr7BAasFs+5I/WJvZIZqBV+lPem/
c5XMUfwq6ZW98v0vqwRxpy46deQ+Iemu6sRvTl1I8CzbhQlf9SBdloRwxhW+CKw5
gODDaOBEn+w9anvixjWvMRmDNNyn4XGAYBCb1fcHbQGtKGtmmY7QEpd0KSq7hQ1C
ru68ZORCfXjDF4ctUvYjfaIQwxHubdp6sM5pIct/FxBzrNYG/g1whUKj6hsKSKy6
4SMm83X1/diB60C1K0W0lsPjhAaIIGBXGiosoWV9IzIIInvaXm567ajy+cZurfxt
vwiGaeG6tGz52NnT7LBk0/XAK1pSu0gBa64EHi4cOWH5uGWSDdZewT6IzXrRhPV8
VyrrnjJgj25/dr+4rnZe8XRCIOjAX/Bi4RTMdIjLADaoWgm8GTgEoKMAgflr1a0A
cFx9LfHhSiXDnyYNj1t18hOluDjdVvTYTWQPkZF7+BrWNKQGT3HZRKigW9kxGXIB
Fo2Y1JrH2BcaJuw1JCSgtNWB7ITIt7B4dJcmuPkI/GNOycgp21U+e1LG7UPBSi74
meZmuzxbpIzQ0M8Cabl/bAifNJ/GMAUEC50ej/CDwqRlVdvwvmDKWNvg4WMChko6
OzG6Ur3hreDtSA4pIv7cHmnVd955lNObDbe90QM4a15U84pkIlC/LG1H1kdCUsFO
4SeUXBUUN0/lL/d8xfWu03Kd1ZyjhaxoMiaDiXMkfFv5KrrNB5lcqXcwxS65KtHw
XvxwaaQuWtv6KiF915/rcIucfj3EakRB2ZGuSaljmWJfx71gv6OoDEXUME9IGaHg
qJY4Z5d82kRzby2qR+aq0PZMCDC+nxout329A4l9EAIKTEHoBR7N+rgsUi4L9zeM
Ux5CNy847KStYt+fXsQQOmv0sFIX+bxS3amIIWNhqyM089RVPq23iNHl2RGSg1yl
LnptILlT6QojsXGfDqqdaYqiQbN/w0mf3qhsGC7sTTk4deT6Q2FEMNBeHgwIj3g0
xiXeaQJU1zgyVWE/JfJcPaZpeYerMOL2eca1OPrZGZ7aK7d7Blt028sV7cqPFTbh
x6Ha5FAcVu9rRJ78k95ULY6BxWA+sphZOfWYOm66NCTkNaUSqOjmW+9pWnIHQx6k
Przt5IZU7KF6sqMUUaNqjdCBXn5XqVpcDlaEC79K8C/d62+ocw/SagaLZfzylt9v
Zir3j6UylI2FnmLdpSIdKNjGBL7+astd0D94exLQkVWasizjFuHNdOJOOcE7i1sB
4BiVw8N5hWkDIdy4ijBUZhsh7L6Lf7NFGsjpJjarmBpeC0ZkYiRqxxJjTsswh0rE
ywAHVklD/wIqXStnqYlwsgGNpNOoTiVErN9UXNowSTjXmbgc26aFojKVsSq7OKuO
Wrxg7pC3jUw6lsKr2nsuPbMc6tTUBAFB3+4FjYFprzX2nYn8klqvSdDfHGI1q9Bb
WWda2R9uf2WBWuKx6Gr02bN36HvsslDRPb4Y4W572PiGQGlsv/p959oyPxauhy3Q
vmgPcdLJDiEE8f3oUF64CjAXpQIWTysuhSKdZa9/Yz8+qCg7jxXKaz4d4WG59WLA
JrPAVPnwCqV3upfkqoizFYb11jg22KKAUMwHVZ1ArQaWA5Kc/UGGKek5gCwz0z0I
/2irBj/HF1yiUDyqEJ4zSoxff1iAntb1cjKEFlkCk0c/XZQcDR35NH7kwRBSle0q
Eatyxli9X3DYVd9arTLydnn4ksBnf15VL1gfhqg6EpJRiaLSz9ZJ+HChZiqXAbKv
2MPJJd9tXdFUDBwK8thth4iPmz+gtze//3/52RN2o2LEw93nuOPRG+hmUIs+Rjnl
eZObUoLVXoZLmXLszOWlB6OiDo+FEQGKrXnkwbTs8IRRXCaRxgk+cww93ohL/yH/
2m5zDENQ3p9Yo46B62DvglIlHkAgVnbvQuSUlSFBvN3THlIGeHSz46nBmYy83Z+g
jJyRqiYdHVbD/TPbOK98KzizdCHK4SVr3YGZniS1Hgb8D/h3kKFOXFxrqA30t4af
GPJwvitNzy++VyLq0qKSVDtny52HEnYqDNFZDYil19IclWR1aL+zzIrYJCHnsI6/
YpmUICpjl6kJUHqW1h1GdonInVOizI8pxwr7dpli2/XZhoWXNCz+IYgULUVv5PnF
/55uhC/1Onqikeeaf97brG5yzDdYfbe40McGB4OcrYQfpBDYqxw8NfWM/sZx2BOT
UNpUWwsCIlDxAGB7jX6o0LiaVNfs6eLLQLx4zEeTnGTCNnvlneZqyhmJoglRUNdR
6KLij/5Z3NNWdFrcK31V87QENjdHbYXL6N1fiW9VRIegnf2MhSvyEDD0y5brTHJF
uDHOLzlBo5makfciOoVgc9d+UqBMLWdD7GV62AkvJrdhyJ9YHQH8ojd5Y9lN9xVJ
fUFL4NTnwqOI8PLpPKnhNziLAYnJdVJsCZAwffStWFIYAHWmXGezlFtv6VfZCIOw
0a6fYe2AFq8KUFjyfOPpZEeyxQB+KUPAMC+5S2oZbFYcX/RcDrVE7lGv+c12Uqpd
Q58dAna0K8ow0qmHOJVy/lUjDWPN6fz71VjdVyLEgusBgEBEIOP4S62u1Tn6R61U
5Cxy+UUuQwhYy0V8sOboVR0vb2v9IadPo4VM5dxGggMCdvlUfO+1gK2vLPPRUOXb
nVnqgsbytMPgcskN+mBRHnzyLeYoW0eKfUNPzal1dulDoVF3G0GQApOanOenQPwH
Zm7gjIkSTwV6Rnz07xoiQFuz7cSaFm96bqyP2cW0YL3Nka3uzmxbfZwq5qsQDRjY
jyb33LzrVsZVxJvnYnafoNWxFuUiCYtROetGIS+tUUTbb/u/bK4y+KQVMKTUzRG5
rKOjA5Fq8KB9EdKtt2tviv1tWVknUFX2kMgWsXdfZeVSCbLmiiLIxlZFsGJRv3Bf
gVoIeUcrFTmH/9AQfMDO7rx5wBmWm2IZoQqPeBnJcpco5qW8hWFRmTDqrM+OxDHB
U2n/4hBQkBrGoFixbVFfr0KoUW7co+U9xIQ+xFLVNC+Z5PuTN3P3W005dVsVqCiy
K4Cd2qet2S9W4c7+nHyuSZGzUPwVlDs7HTIZb2H/daUqV1nYEoRNIXCiT04ZphX2
LVEbeXkB8rhibKY6+hmm/3Jzc+0GgV1Um7gLrTjCfXpDDVvKr/6jPCloupKuuT5P
qXSC7vXPPp4qNnnjw/IwHfeA5xa3g3C/LRvSUgtpo5QL3ehFSffcfJ7xmVzMs90W
311PizK0gdu4yz31o9UqHrStzrDpSidG3mCO+ZYw5YoHUVDA64RdoKUESp+LsY2U
azf83so/kCw2aqYCH6bY7+H1u1JrjGKGbyw68oGVInEIJWrGUor+qSTCn4UIP1ab
XaTjrdYN/ovIQN7ia0eZLn0Hn9SigMcGYOCnIAbyeVOFIg54yI31ceORsfcmCYo1
An+GscsU43kY3waOQZ4QxEFawql4e7zaBU/NRuIm/cZai04X9/W/yWY/7wNTKuMu
fnAwbIHCapRvThmuHEn6M4Q2ISHbaMvC4+Q3PiROrOtsCnIpKlIkjNcIRRpYhBpX
6vGUxHxbkdDvAVhdwmaLRTaYP0RAW8DfHAFc65Ml83sG+CIeimik7AXDzfTBQ24c
8FHcW/gOvTuuBTVsbTYZsw1n62lVuQUaiyuXyovJndlMtP+jwPtWuYDp0xjGECQI
A3++Wq84W+aIZQiIPcir3czt2jLAh3imbhKADNRWleJB/xKHHRZWZWVius18Gwc6
7anQ5WR6cjdfCouh0JtBrCW5vXBOCbSwvIGV58aSi1Oy7hORRJdetiCfj6TKls64
LWLmMDUggUKhFm8Coc7hr440j0dUuzZ96nSryoR0i+BJB+g0iP/FppUlm+rKUpTN
qLiiNKvkB9n4Szs646r8+RNUZIX+ZJUwpFMBfE63wLkfNDY45Pn/5OvTYRKE4RYT
HdaeI8Th/nRRDtYGs+FELpr0uIKfFGKWQk+LLLlV41CdNBjqlxmaxED4+m3Axg0D
smSfqTUNSxt1frkh2XHz3uA0nopj604uWKpX5Y69WlXEs36eO0+272dTQ1P9Tnss
a1h7JI48a80UVk6ozIDATztifJhW5z/nm+CIVlVxz6GWJaqNaPpZhC51nD+WQOkH
NjSj3Jydw+Asq55CQBF0LAFw+XuDqlG+ea7uRkwYgf0XOgb6PYWyxMt1hjJpDoDx
kTU4YnDnoh7/agVGsGsZCMLlz8y9OGhovMr3BgedsdBUsACLMfqQmbMYHXD4FSku
nkTI40QM+UsLGoitFQsMU1TnItyD7mfsyPwhkpYswphN/CdD2u/apWXf4fU+ZZm1
E6J7aciu/R73o+Kb5K6iGqGBU6VMLuc3+0ZjvETshRgEDnrVMVUrrc2dX8vqGIlB
45onpm+bDyavp6jZ08feTul2fHTtoY4BTT4gRx3Q8xaNa5NYOAVnXpHKremLw/Mq
SdkpbW0/1r2Xpj04eqleF6gOX5Ynf+kprqP1WQ7EQ8BUi9Dq+JnO/ZmmPmGPBS3n
csb/D53s+v36x0ClNn9KSJXTY1IhSSFLUaKLA5SBIw5kwrFlFi1pVKMoRS4bi/i2
7UDCPXFt1FVqs6t3xy96+Z29Ak7IYJx6J1pVPxylB6vdRf/l35+0n8Cims532USQ
FXzgNC26wn9EVwbBfFhWYrXjJYiBJ13fRlP0C3+i5Gl/3Fy4ktJRDPQP2EX+Bp07
cVvN6Uk6S1WR2R4nuxXehvIHWHSgd1paH2rtO+/Ct7LeG+tVDHpWECYiHpAXroZH
EhVyEVElUegaJxIAlGXbYo5ivoJHsTBGjKSaBEMfRDW7yTVprVvuOJqnniXmzbCu
rlUcjQKIFHjAzyzHcKpq5sHV0vF8/6qJKANgQKZW52fkZaklPlkDPYm6qYjrDmgj
xx304MhJJJqSW/aOD8n/CCTaT+ULJzzjHy/D6uZYiIkxpXLTA2xlV/qo9E3IYCt6
lpqriIKmut3ag57CrekjDDjQ8FtoqW4pfrVL/FjDbzWfzvMHGra02xiXYvPbAqxv
tQFg5DlRDdRdTWloWjdc7NrdMT71mgj2tjFcpP1DTfen99sIqnFcwZ1dCe0oi8ke
bhbEcjx/6iMcGpoSuCWRvq5HnG2HYn/sz1Glto2+hYjR9lZ8XtAs3cTWX/9fn8z3
Om9oGlzmYiAY7619VLOLezNOrmcIJibgeHIj8lw+6d6ymfBX+bPW8H6XThvSwd6s
IQB6KlvB404B3hYlLTrU/rknFGKVbvfXSZ1QKBeFhZFTK3Cd7KayHp96RHQelspc
l6bFB9UvBh9e7BllJI7eQqUfA64CefV95tocPUFJB6kFMktQ3veBio94sH1ATiGt
PVvapecYkEHgLDxmyJgBcMl4TN13A8RV/YC9TTd353FpksT0qinPdOPgittvxLBk
lAbBlO6D/JXfgkIKMHhgEFFWJVlx1xxl+jYxt+ogdIuMwra0jxMuBamYmTcT24Fi
TIQ2cqLYIcjQyzgCdwCwCSzv9g0axyWvItDz+q6PsO6YeCkFasQe6j0qZoAnauqq
qXfEJG9yJhbaKDil+53BBoYhSQxx/y25QqrEzstdFZ3VQ7P59DutVNlPpGFACr4E
pYbCuHLmYeBkWtX7vSOWpEROnoccoSHDbvilzq66QguU/2V1a5+1+0L034ZJlXXY
WgigIQtZT1wWnarldksW2w/Ezm7GdDG/qnfBDytkVgL9qoJZjkm53rXFbDMubJsW
ZuKAJDqHqH/ed8UMHOB27RKkevEPZbzKNFTBIoCZxWJ1JsURddGHYs+yNNtVL2+f
ZlSb3OKF5MOVdLenESbSkL+8JpygP1ZpQ0UNK1XOlHslF7dIBCPAs3UygTqfXmlP
CH9OOgHCXi+awoISfnnMH8WGVPT2ZQ4mT0sZi9rz9qErqIc7dumngiLDcEK97E/O
WLd7IjPTncfgRs5bjVsp76UBcuSxan9FaW2FpYRRmjkZ9ch6cy9vhhRF62la8Dje
7GpIm2D8NWZDRVFZrX/J9+iSEJxf+yY4sTqnGqo8rL+LvcGi2aIgsBDU0S7R5P72
+BjwLCh6boMFISLGrMfoX2Let4UHL61S8dPGQE4jeTWAholjq8BQVNuvxbdy1Ysf
sqbNuEsaGxPEZyiWzZVP/aEv/iFh4+yRN95FMjLqAyRVZDpoDJYSpZZ2SdMzvyfW
hxalmFa7jYpZrS+tl7LBp9vzNiWT2swcAIArw6f7/93m2PT/GpJV7zv244CjxjEy
DRN8Jp+HzG6V6BVuW+E0/LpEUQzAXcXOCq+Nlaxnch9VkfUYIQkV94RW8HZb55Q8
B8Tas15F3K69GM5EFXnyFZys+FfKoBJ7LLjcI6XYWZOnLzHJLLUPm9mviZMKf/J8
osczocsTf9Wb4a5uu0q3oZeg91C5TeJgtfKlAupMQ1WHFNXVEAK6Nz5926YQcrv1
5+WGpNOwEU4bS3zvraYfA4Ym5gfU1KkAF+jLiaVF7SWTn2zmsf1juj68whttYUOq
OLu57KMftNA5tUlxhNlF40PDuBiQm/eeBBE0xBhat4Vbb/1XBYDsqNQQGppkKAUu
I+Zo0pZP6SPmEhZ0iORWqE+S2Ll1zNSsy84ulbI4HUph2Zr4BswCSgYrurZ7CmQc
/7MHTSCdrOl2KWUQkIMeikKS6TkrTE//IJA/pqB+D7V92Tce9xhR4ifuSoYcadMR
HpC2PDlbZnp+wep1GncS4ZpDMXdMX4b3rBVUfwbtOAa/OlHnWt7ia9n9QQ0foWfj
+aZaq9LLBOEvwMJKTfe78ruM0Kkf8bWXGYnnyptFX3/NFTp7FwzpEnYki+NRIBeQ
V4PvkB0dU0mATg1bGdIeXuDMYLIEZYVs0BNrWJkketqnPK350k/6QaTiJlXuqxug
i6iuQk3ijeNIkzBvcnIeCQ4aC2mC6v61io9t4sS+UIl19AVwfWfbA3LR8Vgc7IuW
PuGNOpQYeTlwAHqwBG9BLK7FXc/7iUwTLJG03V5etAONiLseBJ+/X8JpmFDn2KNn
fY3Z+Y3i6SouEzwqtot8pqRjKCjSJ4+DHrpGSxCqmKthKejZ0GhYZSzmmIdAhO2K
LdAjVM8sekdwqyvm91XLdkk7wiREjoKpHKhBOYY8lPt1MghczAxjMG13IyzM1pv6
KnNsD6oNgSIKwnbseviEsH+tIWWyNwxEFEuoLX9gmjA/gm51QQXEVbckuj+1LZlr
WqQnc2GwgllptHe8YY2xTs+b+QJjc9Fp+PNihvLReidQee83KuRANczgsM+vHwuJ
SQOUETu36sQPcYzvCXZt1G1ZTDS972gxBUo18uQgC4u4KXe4ADMinCYYXfr1jdSq
0wI/6FrOyHwDwaSsMMbm6Fq88l7QSKsKw9BI34NZkCPkA8yLzsysmhwLIomwQWc8
1dujNTBhUQ3ERWGes32y85jK0+qloF+LqwEgVfnteE/avTEGVyeVNtM//2fcXHf3
dhSym0z6JlFC74+SPcYhlB0suB7UOhoTXiZ/ZBRBCM9isw9hPsMDhQnoSItUVwCj
0IqaZoiXX5ZtNmnUMUBmzom3yv71acIjGxotPoPZqBkoeO0lLPreZJOTLA58k4kC
mbznqyu5beRWJNR0kWT0VJ3+RrcZQfNr2kLEfSpvc6sNCZ/AGNZvan+Ae7ooTw27
SdtxZURSWeiCiyIj8P0Gr5RNR1QkY2A10gbARsEXuRf6utz0uPx9zfTIwEA/NEX1
Wy86G/vuNsYxlU1DrLpeuben1s3nzyWsQ7VvqJ3ez7BJbpm7ZQGd8bmsWgkqxtVI
7zXvqhj0OpnzfvMCMqsGL7rF8OaMFUmGUPnBaTHckeayECguJhpaiwf5qSa2OfO1
44ihuRiMqdY32PhyuK3gqum5VfTklsNSg85teJLsJ/vpdePfGd2DOCDcPZn5YdKW
F8EZUTjD+R219+kz++DbVcSGMpZWyjD42MTxCBt7nm4=
`pragma protect end_protected
