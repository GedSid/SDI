// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:38 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
J3HLeYsFgU0SDfpl4LpicyQbNu4rDwjlYVkEokD3iYNk4IVh7IekxZ4ivEZB2l1d
UewCPmfOBluuvOZmp5nj7rer8Ps5zbre5IM37zAbOMxwJ3/l7O+hEDIj6OLCFfih
xUk/CgodxGIp9ypnXmCtO0pfXuASic3b4YEtBgqDOwU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7088)
jh0EKTcqVDVyClW7NWJSj5rFjO9odQu6hZGUOkO+JB321OIEKAh7lfQLHFOF3O3O
pScM0haqKLprpKzsU70GWmgvU23sT8uHvAA2RHw1xSg99sDRBvfKySfRNb9egVMU
Wxi3BwYeC0JAzW9xsiI+E1yw/jktWmAPBB/+4lwhSQNFSn86gNdELIEtogMDoWV/
uZeDfRN3j8+ZXiO29V3ayV8nICr9gC6x0AuqEoZaXkka9Kx52r1OSr+NmIN7rBNU
8Xa3fcdHAYP6gycMT2q1mZb/2bnVORhgEpZHLpYSqmRL54HluLo0VdjLjMgekbkD
yvBaDgFWCPihMoK/ua42RmLuxLhawHrb0AhrcVQluAMEK/CbMtEaLQjUgKOi3I5o
fIaETQGvLNiLvK9BRORKf70/h9sPIXO3vLjBC7NAUP6ER7njtmudfmgtdCQu844M
9vQExP3K1xPyb6Lsl7J4KKMxonbVeIXUHkoHgx5PTVAnIUWkIOKtaG7OZSSi3UCC
YNoJUiz/05kEXKWVBDTAkHM6cZRVTd2ysKq14SWWbBNwDsJTF4qpCX8bmvZPN3Ha
zFhwVq6qrCc5lhoDJT2lC8vNzRsPhQRLiVliBg5umxXDAcRQ+0CkHp8bmNO+m596
YVzkXXMMtF8AYPrJeNHcrAhjgej5I5eFOXSEDho52uwNBiEoJif6Eu2DVNGv65iS
2Y7bUVD62mCxp9Wm0A4VwqHUbzgCdDizmGUk69xqwOXlh4FkJfhK9V1ZlrJYDEXc
UYH2sairCCrgNFqg/fkk8ZxG9EXC/PsWxqQxp6O8I5DbhgSR3+HSX2FLFtXFkZsL
6QrtOszLXkZxljGo6I8XwZ9fbB1zzfsx78DEx/2bwupgZOfEaMAQC6nBLk45G4oe
eOIISNnH+AnI2xerZtsqg6YWlwaowUwMvmwtKqR0dBbxckTmPFJLRpUj3T3R+qrH
/mNItffkrx/cIHwvMCYvvnZIomjp046TdkT2JziAHQgcPVMsmSwoWQNmTG9ihsnH
VGiMYnqGCKxeG5yboEa48RYcMkWyvFZN/9y2Rs8RPdfU+eRrUcYZhG95MU43j3/T
wna+BNhMiCMRAYw16GryLhxJrnP+eaLiWUTHm0wVSa9vgL5pIicRkG0JRu+Ouvl9
JTobcIInrj7vFL0ZT/q6kIY/GwJCoDj7pZvp+BW6+EUGiVxGZ0XsNByBbzKlECRr
T1Qh5b94nRqsFMflnDCJKuGmwud+ShbXGrXeYyuxlGO1JjJMla6Dd4ZPYJVl1qXW
m3846LW7H9aQWuxZRHgrIg8+M3MScjg6iluf5xZJ1H3iiYX07NIGNqKSy0pI6D3X
Yfb1LnyqwOaP89gccUYPIF2tzQ+i2XBqkli7OmLX8TL8xLEXpaKMjHeVBQIdLMx2
c72D27QwrIAGJMGNAojExjoXRdyUSFENUTRS1J6M0FAFCL3LmfCQI/TlvjmI8Vwd
0FNZHOeDHHGNc2re1lW/k7EXaM81nONSVjupM4KN36BVKN2039/q4MOLHrSV1Ohy
l8AH3kd8GsfhizW2phHUqmK9iKtaFwoPAok8tu8VgyTqnB6D3guK2lZDPyKDVJHR
vu4T3OXHlxosYfg5o5xMa8K4W+Z+RhDbwurkpklOHbI2exR05F6VUlvx2252+IFG
UCbuZpG9/onNkZG7BURkIMLWWL9hFqqgk4U/bEQQ8uNFkgZnrGFx5c2CIEGFNjOr
9CJnTX2/WxEhWM7/OmjOUXkIggVu1og8nwZgGZxtlleiDE6Y/uQ+lIKlarf0p1rv
hjtlkIfXH1UxjTu+QCwkeQHREOmH2qpu+vJ/HFiH++68ElFaNhdFXc7NgLhebnL+
nuIwpb1xzm4QkOduncBfZUwnJbgO+j6rMT/i1yGI9U10PtrhfSEOk0GW5giY0Age
x6gcdsUyrEsa3Rz9OZJQdb1luDrfyPFsnuKTfLuPfkR9oRHssFwSnEQFXHEW0jAJ
iYtY70x0rHy9OPpH1TusbaYodx9rDgBOxk9py3y7x96ATVbJ3Cm/0SOCtlMxBpFb
ooU0qa/znnISZGf1kjzfOn+caNkfMdfdLBQ0LUxmbLhuN7SinDkEEvNqeaF4Vi4Z
mz45ZwDs4cPwvvLvH+xmvAJsL1klQnVkyl6SG9mohhOC3HsjVj/r5+v1S4XMA2UK
5gFnLRhJaEw/LGyg3IG8EF5SiF0ECnoE37A8GSdPSB+0f3tTiLoUfG4nHsF49oZ3
AAfBMZ5GiDKBSNT3exrnPNUuwzYqkA5UJwDbpVPhBJmkh3W7JdLCNjHvUh0Huov1
dLPzWaMJgJQe0VTKt7WNJNGqgTK5pKZtuLqP4d+2dyMKTh/EfcdEuNgC/4IACIrz
1biFJUGQnDDRypg7ifCssf4tpezv9ocYugXyLTGuU3U7GFPe49YaJ+5KocQ5Lj7P
smBIf1dXJr3n/kjRY6OHtxXgHot4RpasaWi2ES2/Lj4M2qvTD7mXcyalRf6atVoQ
oKXPSHirlgX/U03y7yFCbIYrdWdA4GrKzhHg56U0Vez3YVpmpmnYuDJB2pxS/oDH
UmW3qXTjK2VqAAsNc4FkbsggTG/Tv3eHC9hJnVsDq6nvDG3XiulfV4+hflhnA93n
LnZJHWJInFJe0sVoRIHatn4Ksw9uBgJUL+uTa3HfOMrSCki4TlpNixTRjZEzj1bE
4K5pXKDhPskQWYR2JhyPnB3LB/KQgjDozs2i2dkPb8iRhBMhTW/hK5cwJz5thCgm
LtvmABuPt8+0PoE7NkE6ijRvbnYoDMtGH4638hr6fc8lS4YwKU6pm9S0W3Rw8ewC
ZgkoaGrrCbjnwUr8d+/3RfRR1/aSOi4Pj5uI1hIfPtrGswct020kA3qp9oVJ1/Gq
iF699F7XLFahpdGyHYxG0YFDmLd1qMbO9fFkkLgcQZie4WAli6OOTGPBQX2kz9Pq
gvMWydoUwMwGd8Eqs/GOKcTGobGTECwMm9EbFN5mw87Wwky+xq3MA0GLpsGufq1D
wE3E33oIddVcu/9+v9SYHdEJeYuXmiu51AtfvTHhb2pPUifRS9MC/jGPSvxzolep
Cw2WCKZ34niIHolAd0FSQ8iWKPksHDWDXC2mI/yEyaGYYLBOnlisuSjWGpDutjf6
oPmXubLtKDBFCUXgNcN5edyn0rPJj2EWx+BlTkeiZUfO5Lu/CdH/mt7Usnaxw9n0
Yt9MeKd/cayLyajZmuoDICMhjR7ptWQ7dKyh8L/mSOA3Vz8GdmHL3fjvIxGr5WMj
zNocS4eRDP4TSLUUydWQMDWHsOvIJXZEZkm3Q0t7B1yFL15MrxFo/EAugdnw9tO1
KgdzFysqh2YnSA7ivIFroCtNrXZPBKc0Srlsttu0ffrlhaMKPeW0jG/bPPFXsW3b
P3Wcg/t1eq6GKwC6FLyxB5hXx5dSBo5JfR08T4fyAtDkaVOB8kRGK5dPVAmv6WnA
nFH4RNeFHkuI7ZZvzh+l+eZLGe+zUBWXdDHhEGAcZ7VktflO2MCvOSjx0rzDifEi
4fnXC0lvBUTBISCXCZsNY/S4V95LfFLme7zkaBCmGOF7KVNplk2Z2r2OX1vhrtWr
sLI+ihyt3i+A+o9I/mQOUs+TaX0YbSIOwuV5Bm9uCiwYAPyl1qstoRKXVnPX8pVE
ez/8GLPTaZfivgdeCUqKGGnfFQElpOJUraGBNcDhrTCfX0waYMTPioh8vshfX46o
d11n6ILGLVycEa0owtNwcHdFV6p3vof3ZrmVYdDz5CgURSCxX94YGbL/I+bkBI2o
5jH5g0FW/ookQZ0syA/vhFJ5ZlWzDFGcIgg6ocn3agP8lkApz8YoZNiqtUwdnufp
RDczfhfZ+wH4h4IWav7UFfYnI5hq0mdM3lG/GfhiI6f5O9xnqe6XDRpegLj3WJX2
Fk7CXlPS99t+Hb0hbeZVhGi8ayjDvf2Xza5I+XCW415JuKPnV98iuQj1GnagVkRC
TwIyqUkdXBh83ZlLzH3wcKE0rVlmQQcpcR519Ib/JvhffhHbPrCoxah722yv33Tw
8aSo0sAOTU1vv2Rgvnf4YKyHTiGRJYnEilMwp+vo7e/sx2Dz+S/4r+e5ihve6yMi
5/FmqwC1oLqB9IY63gVJ92qK0TrKpKHVIXKL3HjgMHAxt2MJbfab9UX1FUOosmVi
Yw+4ujNAY+TXlwz0k4fXIE2m8G5lPnJBkKh/keBvqLBecYCzrTBOliU+gqf2RdRT
hfvc9B3qT9q76y5/UCzdPAc1jczWe7PJLQYj6rEAJm2RL6nmQq+Rl37QEoKbVgW9
fppXvcjMGo8sBHLiatLu8BiuXcPCmW9DkfFc4bEDHCJ/4r+A6sP9buW6r0mWOWwm
jgeuR6V0EIXSdpwmCJoAX3yXXZ1q80gwz95qXrZJ9ru6Bu1fD8/nPD8zCs4pIEIe
zxbLJ7mZQjC4K5jUS0CYRl/Opyu+lDvuQbCkJEW+262DjYICOhMJsG1QYyzXwcBS
d5icNEg9JbBHcD7ut1oIm4g+cGa6n3XKiK4493VmKN8Kc3h8moM1zs/JIcKX5WBr
A2Q78ujVx3K1D5j3RqnQ+oJajgsE/tWt+fKSFMgOwqyoVg0vsWMglMmULM6JJ69u
o3x7YLD+1HOw+i8trI9MhPIu8j0J26NST1byOs2tKZ/4kJhRnoNMD+6U9Q29X0iy
LUVWWb/q1sk+vFcDbkDp9ZZ2Qa3GF/oTyBcyQVY9DY0BE+mV7P9PeHGeT5D6MxVD
+8kP/b/DmU+cR1NeQcM1Ogar06Gp6VwWwN/nEU6PZG/uutLDt/fbNBe73zrNZSUm
Oz0ERc/R1EHkv+P5eQQrPBGV4UiWnTLJ0VXT2ebgx/pUluZw6/Q6GNR3vQQIMwKZ
QhmeN7mk37qbrmmUoLD8tjQEZv8SdjkcT+HqgpCHVhVjcTTJmBku/hR9axq18wzv
lE2oD5tpUv7SN7Adanshnn4cTfc4IbZhN05GCVVR8rb3NwjO6XExsANhqWNPuYJQ
BBt8Rqo/I/0FRuvjVQAIuiMkrIp8E7fmDvsVsoHkKk/QctQTrMYkSRMJlRXYQSxX
rPgmpKaIJ1j/ldgkD94SQ77fyWDCUveBniki/hYcZvT9xv0hdPV2FWiFK7O4P/WW
ewDRHuj+UJM5Dxb3X0xr82/ew5x9UuZ7G6MEt3lSYdXfi9dxSPyA08a44oSp6KcJ
sjl+dq3R4eoAi5wGrNkVxiKiwEMw1OwO4GAtj4Dv0XvqeGOE64t0PJlDcqh6PH1P
Qh32y3a+FmZxoYq0mKzfoOWbA+7MpIZhxZ0roNq3SnGZg5gnYcN/rTBwDuVNnW4I
GvMB6Z4d8N6YNn5Yur/BEF2XexxpF1iDP/zqWML4vIO61qeQdbSNfqkfTzBSen2z
pH/ddlUSTcAZhMGn4axfncgAT/t13e0Se1sbh5AkRLfIR5r3xfn7d95RjmZsoLZ8
o2OFOSwhREx/Tj36yVhUtSQ6fbqTCIK/mK259ayhpuZEpdMg87jEH2xNpvJqKOR4
Q/knUQgndZq5wxaB1VI/gfkdzSk16TYBatbkpw3hmGefzbMvoA4qxKK6l+kraLRf
p5whCetr6X7UNiU391XjthvmUz4mUz62GJKiHZU9sbDKV/BRlBhIxk9eFkWza4HH
Ejki7UgDRQQb/9G3jAjQNAFdhMSeUx+MQP4odgJBP44QGWE55ooD+XkmQgrZmvLm
ImX2JIMe+g2+gkvHl7jcz7+t8mGPcUz9C6IAOPoITaBpFflIR7CiETDwu/ChZGCd
fjUiVGCpeurxLfpt+sDnQd59K/yuyV7IBYAn2UUWOm7zg2l1HIVHEpYTnIGzlR8r
BDyUHMDF8bU11DBw8trjSiHm5HtBGyFoYILGPdmUC7fKsS+J9E4B+G5wRVoHfTrK
QwK9ojpwhT0qXaQrdGE9X0bdEkHrIEHuoQaa290nSmPA2ULwRjbekIo2M0h4U2ih
clzDik+85DuSYpCBirD1/y0/R4hnvmi1mtZ/q/4KWDgIm8MrRTKtQaoJRLee8SoJ
Pfr0BqHHK/aH0y//R2xo7ns8rh6yKg4Bftkj4CFBhB14TAqj/E9N15gi00pI0ccQ
KbBH39Xh1j9DiSKHAsuFDM3pViYl/hMW9snzX74NhdcmHsnprT8KaTbjyJz9Nz6Q
MTQZv+oiAV/8JU4lryggRRfNg9Cd4G3pswypMrLoYeZhbHbaiXV5CIr/uCgtZuWh
O6NTGzYBSxzH834JKQZrHGB/gnRyZD1ghvn1bMVuXpmeA3BATX353AoBdUxGTOnG
ceo83ZwcgAiW5IUwJLoVeKJ6xkJcnoFvOcJwsQtzle2ejHrTzwlBgUjiWakaSdUN
oFTFNQMVHHF3nzmLu2SeFjxGuFdKAYc8tk6RjjesoCh7XrTO5jROKp8x8aRX+phe
uNzoWU/FWMGQI9bDDoWDrGYXzpunl8kkwMQiGpsxc5g7REDy0KJ9MvtbU8HU3SWW
YjzDyLI7WTHP2T9vtJgWH3X2WPktWdeoETGJiCwsWrVQcmEEKccVHRyIoE5N+Ylt
kHc0ceQcfoMAONz9dt4+ZYr3R/2Wd4hSRU5UbTiEzeqcweMYKJd79YhrZUakoTdw
8PoUPJYTLSQUJ51O+XRq8NTMWD+2/mm0+h85B8t5BYABQUQG5KAJTp8IcOQjp+7z
8/1YdYQkHfPbaz+JxWQLyarl3r2n26PzqoWjy6EUMwJsY8FuLFwXVCS25b432gVG
YCtSaj1FosGFiVMldmZiL5Ftl2aW+rzdVgILRyGLtGgL50M8nS/+uP64r5nIEvNb
AQnyIuFBH0TqWuJcv6OK3UL589atAU7/Hj53m6xZOdPZA6H8vgzLrfrtOoFeS5oE
a1RnHvFtfumrNcu2QzFkBd6a/811oCT7eE01R5h5XHMoNd2itd6tTvW/elj8zcAO
gmEGu9IKiBNglw99wAUhFgy2jo3IX2GZf/jJCvA7NlvaXqSihWV8O6GL5rAkUhl4
ZXygLv/1q4oVHwwpEeeB+pQ8ZDuJpMGHu1RQVJwJeky4KQhuds8waXpEsGR5VCFj
EMV8KuCK7xdE2uIZVV7erziaBnDxl3YMJNBLzh239H+cX5QdRi7xZ2I/SHvDw0YH
rAY/DHbY0EHYEb2956YbtIyfSoI1lgymmSIZAky4wR+XTfzdGvgbaFdCfDVlLSyU
4uHxNScNRkNSzh0DAVbpQEfKu2HrGeF/iJyP1jr0uPNl01SKlehwEEbL1EalPeQY
rjMh4OlSD2vqV1BS+UlkecLjFtT1TtY+xXHfQJhBuVsH5f1Sb+/0gts5LWImMX/u
646t0L9Mj5Tq0C+w6mo4hZS0saYJBkfxnhOzn3i5vGIJlgYNNcvff6YN5BH77jJv
u46qY7xfTeYGZeH6uPVC0ZS9W42JVl0InNMeW/sO5qM5i1mWoa0fe+NyZjj6gQz6
Io7ZgISOCY4cvRcfVY4lXnmGP38YjimV3AvAgKs1zBHsoYGFf1VqiBI6hGEQBOBd
WuEFoWBIGlWzcXIRCypSoJPZfN++K1xR9NqDL+FI5JxXJONgXvBSH9D+nLJ61Hrb
p+7q27+7iUvmhJ/ka52+7adBeuV7t39aOxZSKSUQ082rSegRlcjM04T6xvGtKh5e
Uez5kr9pA0VDP8KAGTJdJvFoUueu5MeUORdalamKhWWkaYK2bCSR9gzfC+W01R7I
msrSjKlpA0LUrSaxl1+Rx/UnfcTXSCooEB6nHjdGlwW/9DY64S7lTWOgg3gdzmE/
s7S5gOe7xdZBY8S7Q7L4Kcgy5ZFyQmGtDwuY5/8FNum+EFpLK9T5wMqoQp6OCSa7
8tkhqqb4bybAFkubHSGwhl1fHqZn/87Tlz+NGorhS70QuGe2L14qYU4xoPk3cvJg
Ua8Xz47BwG76YRYrTDBBl6lLjEKQnvwny13yeFDI/Dkr2vegOfj07J+JlXrf3TK5
hWVEacEy8iwo1x2bpiD4MI2MJVupAHQ4jp8AlIxCIh0U4CO+ptBQHumUnVIsQfcw
q7pHMS5MPdIevgdrcgMJ5ZxhuMn7ynMIzkm4vCvW97EJdXwHP8pNYGSmzT07YQaj
EBBgAi8SOsqZl062W+SWu7jHlopjXeOrsvIhQWa5ebU4s95OUpm9RkjXdD0frHxo
j1XHvGsIqhpNsTcA0UYrttnNz1hsAwm0x1NT8eMap4elcNzTU/mSp/hWsYdu2bfy
lj0PDx6d5Byhp25bMvs6igt6J3zS6seelOTjeqq8/i9sJR5vtmC7Aj9T/oNAmAHO
i/G9LFSw6uBNutQOLFMKw2WOYRNkKqtAEuFYR1Mqy2VHQJ6/niDdTaySu3OsA7G5
EjHc1df4yK/jTKEGVHp5AFWAy313/JPeVAwy9LCpheaLZAyGbPkAMbzPv660zaIG
O+M0G9dXM7IDvMJ4ytmxCrTE/3/cKKVFMOBSMsgPcEQFFYAzRJxvMsnrfgiCC/H9
scQf9h1jXlOe83nZk7EcpPLanXRXAAEF7p1CInzAVIsGRTpgHaZkYrGojXqM7MzH
Evxi4N4M3xhdeDck5YaHj0oHDUSsOliCtmYlkqEItDbn0sk2j0niwvgn/7UT3iLv
jJo4O//vUdIZjjUFAqfzIa08I2IoJY1z1VzOW31LqD/Ok+8tRDjW6fkrxrdqqiIB
7Mhf1Efy1K1AzKRKxtVqzFpqL9D3YmLO1s+CHtjsZhWGDA5C2SnoSaYiHFU8JIGY
Or+PvPbGLH8TdtaBIMJec8DzOuQjPhlf5OUf3/DBHRmrDHs41vm/OpvWJsZGEojl
/MhLZa0vMv3wdmSo1ejz+hIvp0u7a2VriCptQ8veBIcst4RwZtF+8w6+a2W7FhhE
huUIX1/fS3/Abl0hHH8yddoiK5CeAwDKHdAFPkCEUtJq9wGh3wrbNuQlPI9TXkZK
WL4Q/EPEOC2KaIL4aQmsqgYUeXWCn712JF967Xu3o5nD6/BNomVsSP10H1gcu3dq
GEW1BceNZOH5T5882c3vAV1I+KMM0mLpDdnr9ftGydj/BJCUicuipUUMfOW3gj2R
b1Mxcxy751ATfLy0WTylWS3SZdO7J0Qy2WKoCGthGe+sRQzwsounPRZhLa1amCQ9
sYGtdPjSJ3Mw0l+y42WvwBbhX8IgtyBHFAxANlrrs5JXWEC71uSicqfiPMYTalkn
gbyKqmbopPtt9Z8mNja73VCQDq/pWPL9rzsb57uuW3N97pA+hdAqiO45pw4tMPz2
YApBs1AZxpOijlk5zmQep+TbNbZxloojkOV1rl4w+FBT7UwbSzONoT1aNMDEfPIe
QTHzMkgyYMVkkTR09m5W7laosXLwtOtbQ11RYXqnfcdH7o4BdzuMnxL/rKuuwemj
NjXVfIEHPxQ7Ijz7HoL6BxTq8ABYMqiTnzZFgwO/oBCiNNJekrM8RFMqrGBoqmgJ
V2oanNP0rxdadMQ84gOyxhnYsLr0WZghQABovvEA6Go=
`pragma protect end_protected
