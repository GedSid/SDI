// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:13 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mvJg6xtnTN3vPdCBDKWs14wz02/ri3dAbZjN6IeauIzcabQVTk1CzkSxDF5tjC7X
PQQLRej0BcmXBZIxUd2xj0mpufrNeTMAVdnZahhuVYdBEB4SrfBj6FhqOANqyY+n
/CO5+HKz34Mr3DZXIwnXkLM6fgTUL5p/+P/rMx4+osc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20528)
cV00/uxtaYanHEOX6UXCIiP4ku0cfUYofmGMM3DJEb300tFhCsVnNZ+NC3Zz8LmE
5cegkAXNTspltDt9vO7R637iQYSTrz35HYQaxMc6v2ufjPvFfJXCe7V8xRxyyq8X
Mi0L515Ip99s1UjRLXhZDDQeb1Cq9zvWMT3Xy3Ub/uFw3rc8t9hkdlLbnYOgdrZk
0vW+84N+fzs/mT0K5tX5CjnrvoD894+T0OlSuUJLk+WzWp9C/I/LZGeaLHcIuqq9
QNLN1eXjvzwWieQnbnvNDncpDEtQ6FkPAD4e1q5spsrg6nFsTvH5fF3CtIbvYNj1
6J1LvogG7Bzz+wEeCGSCTmzmw0v74x6n9yJXf+N4H0F/Gn2mj7/e8HSo+E43TY9n
OzWOMTRdgvUSoi00Tgmw0WnvC2CLIoqkp0uq4l96IJf//VUb0vzh18IOFDfQNLSP
JEdakYHot8BsAKJJhNYt6PBc2Y1eIHsEXRZPXrHz0+6crkBD5mI08ayfJw3Gosft
q5IzXp2BY42oOHS7a0vbgLdypQ1q46HMp7wi87R5W0h5aokIN5BXL8GrTGCwdqYM
Td2ab+UpU50hvWYFA6yeLQ7W3yGlHtFZ8ddz/SrS0Akz5x///YhI4j8EuGLfc1MS
vYqqtj597cS2FMR41k7ZV7n+bONhJzckkBB5cgA5klaL90lsu8aH1wgPehM/GXIc
ldg8/Cd0wfKKCDJRBx1oFhiq3IEfhwg/St49lHt7Q/OYDZEaZ5Q8+yWP7zwg00fx
QA79OSzy15blBpyS6AYPwAa3q+cxJ/In79SbkzZ6h9crSlAotgpYF2Ap2jdhS5P9
cF8df2tdadwBtZ72SJdBqWjLCTLC4iod6gj2Yrev8P2y06yKUR2OzB9Fvo0+8sg5
hLkBVLVpoFVlTbQOYi8FQCUfQZMiOnCvU9qEx6YAUt3RvK6GQ6qjkyouExly3/MW
KeCjW7xAh+O9MphrU94dieAKSzGZXgencOdBe5JLn6p8jGw6vQOUfyjKTDVAyCIt
mOUD6nS4UcYKtTpdyw2lVqUXfq82+U8C7HWo8cse54+lStjk3NJYNDHF6XSKW3sz
msBSDmf1XbUlyF4Fvmys38RXxnf6gdtYr7ucZtTXKMi0vmnYgd3FVL5nH47ftqoT
DqZ1Ts6nElar3OX6cOBX3CWx2tj9lOKTWim9DG3b5cfqKDzbdLuy/eGe7ejdKHii
/OIG2xR/Nmj2nYiGBLHc5bhQHY1ukoMvBh1uG0jBc3eHwefg9U5F4+dFSu7Sh9Fu
Rw4GsBsbdVP9HFScyycatv+fqtIvbV+tWY/JfCcoLS3FIcIC1ux2jcu4uuzpYWLm
1ITNjrrlYBwBKQ0q8J31zaRSJ1OpTvEkOkMMCCYnWiAxMj0F4gcETtRpT9TH+pkC
L5NBSzHFl+DmKiwq7W6zQAgdsC/Kz6LZeQjBEHakRQ9gJK28XDZcMK50aQWLUL7e
bfsdHNtUh4OCthCG4agFMjv0UZDlzgzsfgot0rIrUk1lJRTGvp8xs0/bo8jvXl6g
h0a9+efh6DLleUbGNt4916ZJeWfL6YKkS7qWfCWk111zwoQQReh62xRriXLieKn/
mbykNt1Of1TRJ3e7AThVMdkzZzi1+jMmdPUBTguzcsj3Dcdw/TdXMBGRTCSkPZbr
yC1klj3oINgkBDugfvmrTJ5/PkdmhYTdsTrmEPWNdAuZxUjW11TosvEGtuw/znBT
ShzlpqblEvcots06M6T69xanipw8+QFoqgSUkBTntMpyEi1yr+xTsxGLBVgCPIdO
CnCkkfNj3o2PiZLOM4a5X0zrrpC+f1UTff7VNHfT1Uzgz707gW0FDzyTvyHBAesW
ysX673rWj2Q1Yc0ZF84i7MJ8LHrGQN7NQxDsKUX9hkkbJwV8sMtG4vE8HqY8JDZC
mPuXwMuN3/Kmf4ZY+qn5Fk7nylaRTuBMg9hXKB2x6LVCZWPktrVEzvpVhTdlCPdv
mxA3/oAh821fWYJkIDPJKPyDMA55qHNh2Mz25XL84ekod0ZgImS8KUkCiWOhLix6
0cklJ5djNB4llfbwfmLH6nsbubxjtCZZ3YgPZ61P5mrvKjnUfB1cXchCJMYpKGTY
oqiZdqToaQHyYJxcsDMcxkh6h5ldnEHaup4WIvI74y3h6ZaaCkHOnPLPNkz2dlkk
SsYczSMaVlAEg2KV47/GL/PBT+yGrL/1t3bMXTml4YUa/+SkSQxJUzqV/RiWOcuO
GDa6VmsQ9PS0u0Y2GyT0i0BUtCdP82k5grgcgEcdUAWoZHAdVXmD1QXayTYC4aIQ
nopg0Y7wT5wUp6IZ3r29DftqWLCzq6pjKIZeGvTr4gtxNB1o/fTqkBA9KQw48siW
vBv+97ijppXPGf7b2xQs3nJiODoWvkwVLaacu1bt5ElWrE4X4BsNgZSiYBnPza/N
V0ML1gCHjl3lp2BO1GRJpgCVh+KdQZsSKbmFm8f468APseRh2M6zPEBIX1zuT0+A
60mMBx46Bzoz7aDRgsjbcBHJGn0AGcITvAmz6wa+nFYH7woq/hd/NtpJqHb24FR2
clTK35m9sgOhZ8fTm1Rx8GHw8VK92bDyTOr21eQCCoi+PztRPLfrSVxXAncfJM73
2wM9NaBLKlkALPGzkIenPsmSC3tbhSN7MexeUTHh6UE0QScjJgIIaCxL/3aPEZux
XtbBg6veLegQXUuNe8hIPA1MLgxTGG8Hc1aJWkZyyUgm5z9CBV6sUB2M0xd6O2VO
ZaQcHcgPUJ7F5FrSF1OMLVybvB0QOImh1CoHuVXOLEjhs18juCraD/gtIYlVQO7n
mUaWLQnxJtdNRG5tCEBuk06yCdQWzS7bUztQIG/ypbVahUFck2kpgQw53aoXBugu
5Y60KOCZ2lz63O1QEtF0Z+0eNd79P5VyI9pL7HsI4e2k9TcufHngFQsRjXnWFC9o
H/cvR6xrCKD/lQLJTat11+dCixRW4hONA7bVXWUI3FpfQTfcq+f5apXHuSq3L60Z
zvrx1g6wscg/+j3owrpMNBecZQ1WVevod5QmXBoI/SwgmSp5Dv0etwPtQsJmI1SI
ZXDTAfaPTrcWNb5FUgpkkEUphdUQMIgVCIH7TQK6RwBPY6/9bv+MA64KxLa2ApsM
k/j1iEvxmio1wv4OGN/wGEyBE3fBjZeCacMqWYTmcZ06f2qE6o+RvlaeTUYFRqSv
fSuXb8BirBHm61tEsNDXAkOqO1akIrFxceQYD328x+yw4pTLXUyOUcHv7dAHdlUX
bd9f57llPHlf9fbhsV6C+WDexWTEgMcZZSSt/q0dst5z1iXrxWM2nTSxlC4/ljZL
xlXIhGiVH7I3dks775WXmCBkIKNqAd2cK+AJ0CiVPFRnljFQQNBZFei0Fyhc8yHQ
+zQxMsfTBq2Iqg7eKpcY952ak2fNl2F/VqiWfI3lATGfDwQp+sYk2PgRaKi3MikJ
6G7ieiXqZiQPxBqASqkhGGCKVYDlDRO6kJ/FrIdu3wMjJmgez1g2tVRY8T3WSzjf
/6YpuDuu/99h0hMHkkQ6pz7TkOWKqTF48K8kSRpyEqirBy4Z2YKvZveoDnvWYsO6
VA2ktFCp/jUliBybN9k0t2wCePH+b8cpD0ztGo6cWNfUDll4s9M8mMyy/aB6DBG/
aC+qR8ZpqQv6t2VIbHC07XU/A/emrzk2uLuxq24tXzMM3Rge1qUMiP7sMer7puXn
620yg8kEJEAGJu1tpQzsJJ0t6g5b+UM7YNn/o16wgJnn2Ld5y+eCQHSDYIn8/aZN
25mcYV1sh/jdeq8yciHV87qmjYZvrBqeN/hgjkMu13xFWcJl0szisDiZrWjns20g
+pyMyo6jJe/pCrtG+G/Olx1oJKe6N5hGxMYC0jjOEnN5Lv09JiBDnGH1C1NxNQcz
CO8vumFmGuE03NEBQngQmaX3/X7rDsO+Gsu0Vb+sju2V8azRRaNYIwRx50QIWQjY
7zTO/zhkHN2YHJEuwKD7/vFB1Dco5CrOOdgi85VrUwP/+Ktrzmr8KTeGPKOWJ38T
hAVp/Qa8JX9DAQejeI9FDj9GHhoPOxJI2JpK7vhPgIWgY5fmS0BMZwkEILZDXWcL
sEKloS+E7fUTQWyy/M7EARDzuyE7UxcQul7OYb91vUmTFXsIcIfzjFbF9K++9RDc
1qjW9yBOCrKxY7ab3S3abmMscmofEucuLJtb47QMjRtn8My9dfrpt6Rv+7THltoZ
JlL3AHPElE5yWVIkaor4AbQ0UIOE6gwz4hLuzTzNN9J4kPIix8FPdeQgkTPlGG4C
kyAYh82NoVJYHWpExmYxw0wL48frliO4IPYfP1wOVD7uV3qhwA64uJzIUxTPaVm6
8HSDhfEbgT6GocyMPA5THwAVBhLvCrbSB+eOdRYx7iTo/89i1C/S9Ytk/HtOFU4Z
LHg9wqyIYt2kli+rSA0zr1Ia07rn434iTWF4DzjxPWK/MknvgPA129EF252DRFXT
8cbgTAaOx59T3fBLBZQDxGlxGhBrf0qhrYIRf5kkUjhHUgu4XGm14dbEeKrdT5xn
9/5SLJjmMLwtTazaGPuROIG5WWAD4un1WW0f3UTCcYO1tnA7bd4uaTkgpw9du9Uv
D55jF8Df62DVGodApKearkmJCRo7cVIdqX/3hY87/qUsWYKY3sBtzncmJfG5Oud8
ZvFeWym7U8Of9rN9Nl56ykbBU0H9syLA+ItUpkXXqFuOoLouwYb6L+2eUBj31GcT
fyFveK+txhU3VtBFZp+hAgXI7RIav1vWZYAILmPChYrHVlQLMkxcji7DZIcFsYou
yNp/8U9aq10TibRrQBgcMRtrtANk4NBr69QlKUtEH3n0+lR2h13j/bGjr3iBBQ2D
JnXS1/ot0YWbkjBbvm/+1jaY0QevYr7/5jQkhAH2cH5ObBthcQ/cPqlOwo8+LWrJ
Zgs49lq7IlXnIwbz62Zq5WFDi1mQcdHqrnZ91hz/rLshcVJGilcB3FmArRlZ0tGU
HF09ZF8/cjyQTPbw538dJRwptT4VVQieLM7yb52lk6+usRt7mnPT006ozafD1Aun
MAL6YzrxyqzTPX/iAvZaAaENrAdveK406dbhQdUoU7WOt5oYfn2fxf3+DjnvlTEI
RPLO06xlCpbJipTNog7cq56EHhC+PmYr0GDJ2kikkYslLWJ2Q85dP6OnySIBqdMR
xN091+Kz8cCWDoHiiA2d7PlmmS5W9PuankNIWlqfXmCbhfFinlWcSSAWwd+qMSff
XuVygXyP/lAvHMQHECPO19Kti1BVu7QlzwmENFrB+kmk/9oejvs+wOR1E3eupQg5
0dsYltlFDnzFMteM9bWa4lPUofnaYTILyBSvBjBXwmzAOIZUIhFzq95F6ddWbQ2A
CheERneJckkY9BPU+cGPdSp0Y3mMDpp9ABsiTI/XbsxeWltL8FypSCWu7cmDzK83
q1GLGfWCRey91vwj3luAR8Z8LVff4p3KvZnhPypyybtYsis9E7eSvKlZEAJG+DHW
XntpdgsR2nV1C3PgMP7Qr/3AmT68woCGd41EM+UZpVcSqhMy/S/lBm6ANDRsqh1U
jEF4IBtSK9BW7FOUG95sNytO/mx6hIcdXqy7CqrO6oHLgYGXjb89jYXiWSpR4way
3xVfGZP8H8iecFbviXDLp/O6w3D2bLdbTwCH1JeMuQ6rFYEVcWePgjUe+fOzgjjj
7069Qj0A7G29TTuY/PSoVjGJSDALs8sfbCK1IfMD4OOPUjIkBAKEg3BDbAcmnKt4
eTvVjXhs7cRqp8bRk+eaobQ0hzpatMzrCrFm3UxYCZdARUccmN/5EzQBJwCOv8FF
9jpNNyA1MDe6lt7f+mGGCalIUBjUDrIAYPcQphOwnCSjT7kb8tVXrJUPXcEeh72+
nGnx1oMX3CQqsO4MwlByzf4FUFz1aKkvOB466/8rqbuiA/JK39YdjHVlASAaSmbv
VfgfXJysvOJwYe+ikVUdhvnOESFCaBVQtqpX24ENqVKvOdTWRZ9Zi+QB7d6jwLIn
MJoE4cky9l5kdZLSoRaFsoDh7XR1U2jOezvdWKVHbZ1QrQyAN5F0bJN19hfonnZL
8iD/eTkcUD+z7+tOvzU06oioijEXwBnRrbxH91lbVuCVZh+nPnSnu+9NBoqtL/6l
/MiXd+j/4TG4pKOktefse+QAybZMhlyxJXLBHUx6rJE/5eSPvna81hGMONh6lnc8
UWxBhAHC3LNJjIldD3xQD947gjMCgYJWS9t/6RXB85SIQO98WAQYuD8vAsg8j7p+
5TYQNaAlvgsDsBPUXJv622Xz2IOMov/E2wVK1gu9zOMOwC7LhVzD1KfWroj4dPbm
wOwvccO3PFqTKz/PJxdH972hCL9Qmf/VoaQzhUBjv0iHMYmpObpSvZ0Z5fhNKKzu
BKkfQergpwJhNQ0DyI7I7x7xqHwnK1/bF/4EwOQlAtwLc6QJE9XZEbptAGrGrGKl
SZb78j+RMrrt4Omw1HNY6vh5z7Qy3LAVZi+5fqpN74kl+MLeDdP2SPbgwVh+07kB
TPrrkLuwSqSOwlN8zPmAE+47xHQFVve59IBKPh8tmPV5KKoMoGOWRoHSy8zoykTN
Bib5sS0mBxfxC44Y0Mowan+zB6yvywhLqhoIQuX2NNPax9ykZ49g2tUf/nEk2raz
MZcJP/PaBVD8RfTESHHjFA1cs8EdqhLeiJ3nZE8DZxjmQbWsRCL/S1Gar4qG0Bs1
BD5PvM5JKOwYmAeUIQAA5LLWxFeeZ2sAhNio5R5xXw4+GUU8z3KuQiTKmjK/Cwrm
/ycKafpPer8i/z6kjz9+TOx11JRjAXAjIQl9BKkgC8NCWVZ/xq+W/WG3Et3D9loj
PNtU5+cgDGADDvTBTW4AGnJhqS0VFG0bZSIRCvdc11FsoHovEcUcbbUsVuyLIZSE
/+iKMWGULr1EGJ9j2YNsvhIEctNtTjQRjyfeHSzEQ3jInOdPNJtW0G1qFfQiSYnB
uxKft/9xZRAbdJZqHtzkfD0xGo/mQ/qsk++5y2zTeITsQ00DsiIzZQrSeCf2De1v
WBHw4IxQqWbfPvfHx+nELxAmdAZ18XDRPUXpt4DunI8AyswWfs3SFjOyBwitmbJb
VTRecLQ6OC2Yk34Y49gsvu06BbQNqI9W4L1yqLOrlHeUCfGvyNLghzt+ydt39pYo
y/3HfyrpaAdE3j/Phld1j+9WVzobyoBXVmxPlVn8dMYPdAzUfHkKOhgDSLH8hU3K
TFKs8g7UF/BYPKBC6PvKtSTf4pTZNGrmoD43gdTtJnbxg5jfSslbXrTAPrKdpG6q
K0I+MF/JjJoYecZ8M53LQpxkT9AkldZBEBKnXEukMgkoU4mXj2CBZJYffx1/ywTF
w480TKP/8TWXFSakJsHGR82qVrjPXtws7ZH8JCobyjKgZ9plk/ld/R7hPAsSwxVN
o+vgzf9tXofOEVp2qRIrX45b1G89ZsGQ0MZBMOc8AGXmG52cbVVPzzGcFZ/bHP55
Y0QhQ/mrcswDGcaRtTDb7FLzZJTMDJ9nY7GpNNq7+grEPSA9AiiCq1eN1cjbiGe+
bZ3sTcObkXRZeiJ1kPVMuDIG1Xt1b0s3/4tcMzQJIs03fbuI1VDyCpd3bGLAtrrQ
bNrHRR33lMEYhLHt/wm5v2uY4YtT8Kn7rrkRPWK0Eh5ZtbYRX/CbkFJXodis7tV1
6KAhswv68KRdI56/KjLvLDZmtGGH0uEe2OYQrmre+IEzF9/eQB/ytGFSjR1BAMN4
CEpz2peh41Rawcpls8MgE/WvWeB8iEWqKqrLhcL7zkk7Sw6JvhBNM1nxfpJCpIjn
c7Xa5pq8drDY2aLlpVfg9192xOdbTeDdnqQv0TiDJlwN/XJ3uwtat0P1EGqpGxFY
BAd4rc+fuHDfa3c2DM8PSLrLpVHU26ojTG2eNgs7VbE0WRYR3ciD71VrBy1msGc5
HKP9iuhEoJu5/64j8APMgCSXtC8PpjYHyt+dEaekLSpcoaTAvFdKTHclgrjTg5d1
lbFJreUoTlxg1tAWAPsTSzAv2dtDiQvBdZ4jog16fNmWR4oZ7G/pM37MpZUrD4YT
IS6H+OFryOKV9ceUPl2WAzqe3x8LXLYa3T2qq5moThdb7nfthu5jLllhrihN37Uy
QX99xisLu2lDqWA378/Gd3y1AdgSWAd3a+LXMf2dRfEq8//amgv+ZYSEgU7Rg3Sm
WKY06Zz8Qc1pHfs38+K0xFrGfaGFtJQP1NN0WjMhpU0EtYQNgZBY3+AWnKPzCXqP
DwcKUvlz7kks/8vn8pvU6XoeZgwPtDM+1lgefEGlKgR4AXQ8mWW/gqzvlAMb08fz
KNzrdQs8BzuiEHGgd7IxanjnJjYAkDiY8zij6hMZsxn+l9FPGQiIoDdgFlGqNw0r
EMfuDeG6w+Xkgfi2uWrq8Y4lVeFei2eazTUpTt6sDaPe8ZLKckFZEtWP42V0rGlV
G43JrDpImlscTAK5BpQWiymIhaoELjvzNNjg3E6LBBiTx/UvOn9w6GRgPcr6wGzR
YcjYsepvVzeQkO+awL46m/qswZVqnt5vy/H35x4a7ncWx38hIfOnY5k2NdhuOtSq
jJsq0oUqQYzNFoikJXksvf9+6VXY/DDPFOb/qayvi9bqSW8ZWpDuTR2wEwBpEiNU
wEcZtszMLkn5SFP3FvJCnw1H9WaYdXN8Cxcv3LjNcReQlGUiNP+DYGL8u+Qam0jJ
JXR0ubHB0YxgznycstRdvkIQFWeH3o5ZxJkGsydSkffJWer4m2jY8ex+2uTrEZ0R
W22nm94kcNSiY8qzIxUhi+4blpjn+3BAzPv+33azNaayQcD6bHOnJ0zxkmAvtnao
/BG/uKHBhnRai/kjFwDSNoHqnMvUOwEhKvHcL/+8nmsgkGfFgEoU6chY1z6wgYm6
TTyrIOIzF/BASHBiFDS4AzdFrSlfxyXAxgH1BaIFuXzeSeU2rKuz9UKSTaP57rs8
aM4P0roK28yNUvykEqBSKMX26/uBB8O5dmqudmfWsenXmr+ZwShJu+qWp+t2uCKb
G5uFgg6z5Od9EiTVbcZVQwVIaTpoks6DW2Jw8K6ONXPC3AMo1LiISW2SbhWdwY+/
r08E1McQWYGM3iODdzh394kyQdl3UWPE7wGAM83VWG0D7+MhHtahtiBv6w7AYABm
X1XbYL2mhY8lZmbnolUAJEQOQEVCo+4Vp32LFioicMSQ+Tu7QdIsVpaaUoefpcOj
7q959iL8WvKpFtXMFZ8GIQIB3G0HAt3ePh7vl5JnjiEQipIgW7csFrzwHQD2NIWp
JjixCrF2rCPloJNb8eC6aZWOORIssK6FwZ4V+t+3GA6gJS8/4xllqVhcy3xB//g+
yWzNzSiaQXgdA/OZdefyq6Uc0Oyptlc2X7qEutQpO4qFHl9tqXjvnDJ1kCevsfQV
yrHKs78pXTCpP7VWcils+J9Glm9O7N//xy4skmqLCmPKd4fvlml4ixNP+ei8RDt7
u6EUXsmKd818bKepFPzVQcMtD180IB6CtlXhhAtfLykYbT8ceW18O4I2TU5aHb3Q
7J52DsGs8BCEhGRPOz0wOtKt3YNjNVs5sz8dbyjSrFv9BcNZqT0TJfqLuvg8TJ6E
+yJpMeaEMC01hjtYupxHkdV7a4g4VxVlLFYvu5dkbK6BIkwMwR4a4MmrobSWfp5v
SYneaHLi0AIiPNxg3+2Isboab+lCYzJLJKCr/J5GB65xO3I32WqgF+FjHJQNSb38
zaLjwf2LnMS9EJH266eVTpilHPCe+b18D3IyNUsSsYwRsGRKlbA3cCyOZnCeKwzO
RG8Yut8bALJ6eghbT2KyI9AsCIUYlDdEaUbNvfE/TgvTYpk9mA30akAgyesXnfvR
FJWDTCKRVcnyzzv7WDGRp6kNInqsGgo564jqySQgZa5Z6WACFHixs9IdGeO4kGiP
l3fcu9qlsNYc/jxI8VDdrtZcbVS4CcmbZTTfb/+lVhwXF4I50SCJMhIbDw5zX85G
Ml/M0UbVyPZAKJI+hNWSULN9m4fvL5GSlyF/sayNhikW8aNTK4ExLVzk2vSqOb8J
XmMdn/Dt1/489tP3AgoBISsa08sTzFun5+b5mC+4Ow0BLEcuGOp0KzK4N8+rIbzo
N7mqqoukYWqk8FcgdzlN/IWV7n30CS0uUlg7cAndGCfIAd2Ym8QsmrLxkd9r89d1
hBDjT+tWwPAX+tGjldDllJUurjLzMo7opro252HjfAbl2YYzTQ0dQWkG+EiuZvfl
fWJsgv9xMDv8+rw8Wq0WfhwSpmKAdJbqHdLmuhnutL2M0cDSBi1wpjLBWCTFt6tV
Pl+SMbxV/ixSW2cnrAXlJtoVMpHGaMUTRJ4XjD6oBcxM0hdX7456fo5S6m16k/v6
cf+3wmWdceYkEQlfS2NroLb2i8DIBOEohXVwAX84PCcFC686BV29daLPxJOyt3Aj
pLCsGIUJC0iMy73/tM7iBJgvvN+TtEWpwDQsZ3S84CnRIQ+yzj7hHwcxGHgiyUIe
p3xx+Qp/+9y+42Jx8gKXsK9/mTJ97Awj9OWMjj3sYxbY+Dav2QGZhGaKtW1GFoTE
60AZyqZkeQ/8rxU69K5ep29RXO8fyW5/RpIHRlUODsISGHqVxtDs1OD+ibhk3M3a
ajvp1N38mSU3569m04OnNtPiud6SVf0x/er+ye8VAL5KIhOt10JaF7WhLlk/MINw
1fogvCoLdp7veMH0U8pbRxZ9FEKW23LM9d7Y8Jqe4SQKKcrJ5ppfuwrjoDeYgWkQ
OXYeEN3YtlIUzlQ8LvtF8pWTmMJq9aI/cbxs5exrjgbsgAmDih9ta0LfUrdqQ6bh
Qr2EIJRJ/sV3zICK3b4yoosx31IKt8DtGRR2m4NFipYkjXyVU87udwoma0yGgqcp
wfbSVn1SXh6VQMYfLhuhJfswTV4wdquK3Rb36m7Nb3cpkY7MpK+jhoaoGHiTYYKG
v5rk/2YdeZOUzi5uunURAZF2g1qwUfxKuqKmYUCCEcH7jcTrHmYos/mpIEKt+dzn
enJ6Y01C3hJqzjDall88LAXVmyx6QyFJfU6bE2f0KpSKYBqXIHsvMUkyQhHJMVVo
Pxv7DV11LFCvyOFL/cn+sWpZvxG2rrj9IYWxK0jyazX9YgWwFf7ImBEz99km+oU8
yxOZ9TRM0YdE+ij8Xqe/zs12CjgpOYJMkSitewyTdtlspZaFltDgxZQO17jmJXYU
xVBjkcj0n+JctTEBQ0lle3LxLDA8/ufq0RZ8sdc0+9KMtFc2rJjnAXkz34Xic6zT
vu0+nqxbD0NcAW3pjJH5IH3ABW1S7HEcUvFIkCiN3Mua2KUPOSj9D5KelVqV1YSQ
amNCmu1DizS4UO2xDZabWatm6RHRWp3qd31gsJ9A5AX5gvBjDOKaDEK6gNCR3BBg
95EN08vi0yI1LodZL5KraRvNYxkLiJj+gYqMDWvMJ6x8RtupqMg/7UaVx/1TSTd+
D159QblwehfqI5buP3Hs1VPQbet9Sc8zSUTDlT7vAUW9Mjn+G0gkbjjOG3x8JsQX
zLL+20+Z2DxY7TMM4pKTihY/aM2v0VyIZ1qcCwAuYULgaQAyGkll8n8CNb+EDbF7
tLEYWDCE+VA5qMaq7SmSLuaGFin651rfZ5KqlreaYnphHWg21A615/Ky94YSBisp
xVAiYKP1qyJb6SaycPm6LZU0CmsZ1hFXz7UPxGdFDs99lw5tdYqP+ddMz3G+Q51s
WwXeRP2bnktElSuq4Elx2dg++3enObKemlAv2Zh0y+wJAdeo2KU41MgQoU5vmQPg
28n7+8Mj3/x7umGHNdi7PMuycTGZjnSjzcgRNHeRCCA9HEW2JV7K3lZiAGcIC4/R
7aX8IHzVDmjtKsl8z0uFrM1aDwST96aDsUtVQU0er/7qnigNa0X994JmNzOnCi8P
kIMYSmJrI0NVdnFBjacpuUFEFUtwWioMYMn2dCrq8G3Ew2X/ndNAGKpMXIrmgCpo
8v/H7xqz63Piw9aRND+O+OfPzyMXD/01eeGvXp9ygeMAzNAsKD+nxj9jOivzaP/p
yYRJjbHzASIllkj/nQ5GsDEPezxkvqeLhmDO39wY10cyzf7u9Opx1+IjmOBdKlD4
NHczz3jpoS5VMUjQGKWEi+82eR03Ly7KLY/gYdpy/PPdHjcjj7ENIS1odWZ++A7u
U/eKm3TBH9zk1p+88ReJu6N+tbuA9N19n/UH2sETZOajoL6hfKJMpNle86tylJz+
y8Kdc4V3hN4x5lngXv/r4FzBWmEJlo3jylqEtKSbClErvKQon51pjSR8jmtlnzYS
mD4MuzemXMwpq80HDAhYiWT6U46ZjUOOrqi9ndaQI3k7LM71dVxjNPFDdbg9vch3
BdoDt2Hlm3rqU9AXDnEY4JNuo/viTpgkjoF4cvXRl0oxYgjzEovnQo95qdvAGmkp
SxTp5JlFgj0z6g65Nrl7lg6ryoJ4jZbFTAJzo57pnbR68KDatfmy4vAqaiEemSb1
SjLHfit5apBRqtTwEO8s8awod60TM8IaCx7rMuvadX/D5q54JPdd0lsHA9qF1hF5
ahCy0gdI5R/UrBntefzgZm9Rh9k+yjVINrV7NgHc7CN67bMvNwkz/o1Ijg06CLnS
hhdPob284kVADwt455+ZlLyL/0Rhit0jsdF89T9WIVtFN3+g7MKpEHZf7MzaDn46
LeyCxO6/OcUK672ViRDFe+NGRWje74IG9bH8eQrozpg8I4sP213tevTd2HgtUtbK
ulQDTBUbCB5/tUaZqpfolBWYpvigAWJU0wXHr9spcqxe7Hb5Ln7CWK5jpJ09RE3H
oakK4DbpMxyoOuAQsx+ob/JtK+W0w209sYAY4MophQDQRmeQc+/bwaxriIJxfH50
vTzw2BuwIZxE+JLpti3CzW1xIVRDRLPiXY1EFW16wCZfwJd38WiApVjxBe36JRG5
6mrdCCiC0Fwrsf57GA+uznvidhlaOoZvtoiYui6EmW/X1tm5CSDKsoTRmvcLz5WZ
Y5jQgyNXYPj9cJNVK1/EwWVSIPsdiiuehmc9b6zzg0WAFavTl4lwcpldYqjUqwEm
3SnBPamDHvGIri5lV92whKayFpykE4qi+mpWnQ0aRAxCeOH1nE5hi0z7faMJlmcd
tuqFgpzAawJWejEX9HHNmJsNZbHWPHi2Hd4Y318Cu6b7WBVVWG5zicUv/trw9K2t
i0QesWniG90Izp/KsJMFv1mCVurTz4p8y4fWrrvfnQNaYgGfV45cJB1zmCuODFtV
XglkqtBXGYIPOz5eu2m1zBh0UiPSz4M+WKoIToyPN8pg7NzhMgM1bdgrpP3idS/N
eTpypkN7Y7q03rYCCH7gNQvCMhPHPbCy4VXWEyquYui6VfbEFd1TIN2kvYSJyO38
gXhYVlbcRUnHAn9L1u0tzk2rqUD317SmPsTsoFiZEm3YglawXqi5SOWX/2Jai2Sw
A6akqC8lXCXTZEROM9QySHhrTOrNGiPVpEcbO/fScOrpmVaA7NlvHBYqQnyPMbqN
mChVj6MsUWbH4YA+IW+8w5s66Q8vkxRkcmzqLGVg9lKlQDSQ9VqE81xtshoznAdK
Rm3j6jBJSbtaKD1t3eEwXhEovy8+VriALgkX/IF5k2Pex34+Emd2hCne0QWy6idV
TWaH30u5pM747oEkfHpY+ekr+kjIgOLBU8rK/ejejdF3MR3eT9V8UPH39OxRA3CO
hrxrB8X+yG3Xenh2zgScVHkaPhSPXBPr9HScgYMuUPt44FuILnDPdovHfzL+BkS0
Nsuvangmh8OoYEaXUJU42yntnb1n/m9Yd7qfFHa888dTx0TPctCcev96gdUh5PXq
AhYxUT3JN3drF0m/pn85u0FI06Pj5DwYUhVh3auS8E+r1saitBP0Yn0A6bL9W1N5
f0rfUsZgQGo+Apu6eLoOjosVSzUNfwOdbeF6v2EDSxm+7L+aHMODYDP4TI+hah/Q
cmkL59AduagIs23xB4m40uzIRAtSsg4qzeEtxM0jycCD1GpY1HsafZWxIaCXjoBI
glAjqJpWH0X0eMeOl+8K+jciZlvVKrXqzhTeT9PZwdt0LOblH2spdDjYR26PK6kb
ex3uAuE/DPZViJhFSRllNxcEKmNp7aItYC4YQ22qSTyZeYCKAVkYR+0oJiHSdzvf
j97VDQCvyWvxMrWtzMbcdR29EALjrL2WfnJ6e3tYHQx0zPDqlOR7odl8krTpxbgt
nL439FXidPMP/Gmd71SEra5EBzU2pyyT3EDuVdPI17raZWJoQw5lHig/2Ax0KRFt
6hAyhc7lc+d9D9bsE33ftOweLPF02sKwIz50NI7Z3q+A7qarH3X4Lf/8GAv1iehT
rLvD4x+SdbTd6m9YO7oiis7lBkfEZRSPRo0X9CQDg4JF1u2xo7xryZCnzzgIXK5l
DzQvF/j4FutqRKHxuXFNb8V7HWCRgXTBTfc5GKCTVFUUbm2MJ0USRthqPvOV/lZs
82Sx7Gtaw3bXD899kfVAkpQsPOQvQRbgaPI3pZYp1N8IEaDq4pjL6pUZ7nP/OHAE
6f55Qx39J9tF/V5ndt3X7op990EAV4umTJBvbrOSCUAXDPUFolZv7Zzsr7b8HJVF
xYAKqbMNm+/JSdL/Xni+hUFLBJ19ekC5ttFAvZpmRoUKSgSlFjSAnTBB4BGhVyc6
WqOEJcoYfQ1ojsu9UtHZdcN10fYMsLqpvs/Lbh7iYWb/AGDmw50IT1n5I9xjh3CF
dWmwFKIwkRBSjBXuypVMc+tFxeJyXr1VFLe/RRcYlKdrnfXMTsuZmL4n15MkU5l2
E6Rq36Qz1zqhGGuxVoDX4+10FZalNSO6mVaB8rnEtUtXAhoGaQLTbe6S7eLzNNCA
N1fYJaCy66UKJzb3hDXHEZ5KdqlxLJ5y+KdU3yHpIIHIPOOiBvuWNW/b2h1H40bU
U1cMbPsZfX1A1fcGPhkCObdvJ3Aw0RgB2q5VvfFMcbeq4PWYWIGhIEp9nWP3gQGT
Rd7JRZr68zW0j7bLPOO7iSMcwVPfskNkqcWHPneCPPSqnwOedqBNOyKWbQVEvUGN
/zqK7heCFDVWccpCPiaA6lTgiKnA3Ja+AE0mHUMeg81a7Y8ZjVLSGU6Sh19HS7PT
v0qns67qj0Sjsxy+GYJsGcdw4PgN2DlnaPe8Qg05U9QeQGLo1A0UfwbCaUQPqnJY
n3PJVDX9p8Rin8nvoTblrkjDdpb0XyNo5zg5atn+JS8yQUneh0PeoXAqWUfxByz5
a1UDH3eAdR15i73bNIRvH1xQXhpUt+qKw0Sr7FrMwBvJf+w5iTADs/jOWTC9ROvY
3sPomD4OmnXi6G5mOgrhArHCcTrbWJHFJRCdQP3pUFuJCOe78LGr1Ysz078OxhNS
QD6VXhXjhKDPYaG7yX63/xw3bFwa0WftI3a/WmlXrOiZKPy3H/O6JwURSfGyqjmL
X9AjXS82L4qL5p6tL3K9MhJqrjfMpI4sE8tmSk2b6F3Sbmy9u1cOBM2TlKPTZyZX
os2bgB4MCZCmhqobdImyxKG4qBZqzEDmA8aytzLOObbMwb2/WtNw0xGoF+jhLTsY
PjpuIdRj0bG7ftFgaeasXfLYaUoi4pI/b9Ukf/k6EkNlPXz3HZ72VgwqxpNDoWCH
7mcUZjBfhPvwv0rH5ryHVkL3+5hhvNz0Y6FRIFudNf30zteMN+7zx+y0lISyKK8T
5zaPZDXOuaGH0r7vceHaI0YBpXLV/u1B43rknCizWrAR2GInCmrZ37jWTAGG69hm
JibkMEB5Eq468NBBNO9qBgU7M5O1S0Ke+WOSDUtJ+SuBBPjIREtLFEXO+KWYqIsz
QiwSf+d4GBMt6FjSiondgVFU9oIf49LkMfWDz3Wg/VN8DnhXC7qEAq7caqnvczTe
owYbuoi7Ruv7+lvP4s8imVexNzjfXio9oasVQBEqv+XkhhtxtcbJBb2pnFWOU32M
WJ5mnEx6LPjlRzh16Nwh30K9sLAlvnO/cDivpcPemCTNo4/KrHsRkoN7xi80wVAU
F6aE3rtLVyhJnOtXhoKDgdqMFX4XbhylYFukVK/Qy7ZHgropGYtF5at3xCMf8C5n
wlNPO+MqSXtzSUNIWxDPnHxDRtEMLNOXlChqfCoJAjwUNuzs5kDM+EwZeDn1/MX6
0Jb5LMQ3qsgAKrrQpc/lkfsuCSHjaqJ5E5mbFyPxuU6noY3GYK8Aj9eCbNvAKgpG
WsDGMKMMIjVOkkGtoTDLA6RTVyzykulZafr/9wD6690MSL+HTHD4gevjedYLNvhl
qr6ZZApHP27DIKG4MYKXXBMTy9ns+VqpvKlKTcJpfvdKDhEuB3kQq5Yq76wvV/4K
prHt34VliOUjblSygzdZZIHiMjwrB+306hI8zL7/lD1sE2vNRl/0SMrlIkfwIxpz
i07aK/4J4E62LKDx5Xmp6/hMt3iHsXKN7GgiyRBpjly7V/ksnpysQNiuxoRdJRJx
qq8CSxYC/+CCaw6Bx+eDOVbqLBOE8Z7k08UcIyw+cJpTq6hlVKDsJwa0CzskRQgm
h6+V7N+j8fj2YEhloyh4+B5mH9Own4/OzkEtXraewM1K3N3RWQmdENAtsNTJ/dtp
qhcHlxyBziFdmALIU1Y51TIdnAy7GfnKrGWkcMK8mwEVSmAwlNE1hux9CFLhvatp
RMR4J5b/p6Wa5itRxnuENVO0Ihguzc2JPaUZIVQfadpodvvTnUH8e1bhh+PQPcp0
FGv76GJLANUus8x1D0d2xUq6jdvBnvQYCCIU4azkfcvjL8RaGGA9TpDBV4bFmmwD
hHsTmuD0XaH9gt7vbA3zCpHrPB11Y+PieCv22n5OA5yZT+Z3OSWYXrfGwl6Gb9Bs
xLGtTPe/28F7i3UGnAiEC4AhwF+5H3yBJWL8CIecub+o/R3n6AvoUacKnGMGag7Y
dRHQhrW9woSHN5yr2T4HK4VEWBkCkjkdiLczU9exnkykNdn6nwSk75smDzs2OeOg
C5Pndvpbla7kxouJ5E8lPlBE7TNwhV+ZeITEtweTPQ6isYiy+r61wOa7DkSQVAd9
7fyhLP+RgkGAU5wAU2IlJh+dv1RfgrkOwu0SF1PnXRQf4vmlGUtEGA54nObvGhzS
U+lHR2ILScs48fvhcwcLwd9Mw9jsVA34fhSrNj2jv6wo3zqzLhCsNqd8eK3P3vz7
smZ9yRNjDE6+LBHTQmDXHrhmNucWK7jGgryXLtrnFsrObKbY1GAtpwthHeCBhEw+
yYt3FhSS9YO6UB1gj3lZCv78YJa6+vq36pk11IaimaZyu2zCtGeyv9YfkzVyA8aH
Q/tasFTXevBjl9V5QQV5OcAMfsTD8llcphwWHT0pj853E2vocCewNtovOlHRS/EV
tyO8TCbsJanjP4lEQUGcvlJdEtofR8OpqGqnYhoxzI0fJFWcY6WnZCbCDeEx7oFX
g8k3sJbvArttdlnyhfmE1L7bAaVD8Zr6ET1Fvc9tHXHAHjhruJwzDycthRL8hoQS
FzZ9cMJnFNHS+VZ+AuTa5RHeXxH0PQL4aiF2knEEAvjdv5IG81LtSuMeq8brLTF+
/zfVwy2384/cNP5p4VyV0lpiKUJvHas3prui+p2N28hyowmF53Ey7cyez2wuSSfJ
y+E+mgcQFLqO1v5u+opp8zLrIAqk+a0dkume5tlk4O44sL82MHvGDQ7dGxUru5th
un5seNi8pEvpNZlqi3278EC5zbX/z1K0MztFBC6z+XBJiLMm4t3hYD1Ym1UIy+/I
rWMtK/z9VPrqk5U/5AGPObCHQSIH239R+fdpJdmu5p2Eg9naWGK6hL6JAQOPfhpI
F2HxKzKUKCYLnEV8sQ8TPSs55qfgEwg/S5k7rxa6G8TFdwSGzjMlnRNxwvmYP66k
i0m2iQ7mS1bc7XhufxxTJ9QRFbFFpgr9JcA2e53kA07bhjv2kLP6b+sAGU1bJ/NW
mAaoRSLHIRrp3dFKHezAFnl4mGP3DKjQPhJHaWLVqNuOah+Bh9lkzbCTpUKuzdZI
qHluzkyzNGFLos5l/JhtIDuZBePIrz4wnXAM2/iUhW19lje0dRt+gShPynvP9576
9zJ+Ryi6hlML19Qfr2vP6XPDdMDBEPJjXHkq5VTIAucsS+zT1iKlHAyaTtR8U15a
LKuWZDbBYGwE/3p6UkL+z0PqYtMuREyV+W5On+qukimroUeGjyI90pa7v/e0joQz
dFlC+foKTNv8KiBdtJVTeXPb9SD5B0AIMu+iKSoBdItP372J5uyfDDhTZaS7Hf8z
brsysH59xU7pq2OPkQKupOBxnyXFrzFHY4c9h28DTTyZleccsddHGIsZRFPyd8Ug
2FjCEW/jLvo9YZkUbZIByyiGUoThx+n91zZu01uNTxxUcE68ScTBvD2K4MeFV1St
BAukxyECULLcDXUfi9RBAdtOmMHwBohtrvfQPlZgaffHkTQDyfJpVJkg8ewj2ng7
jVGqbABaNQz4CSGywMzsJgbXtSahx2HiF3XDq1oHvzdXqaaYWpcY45Ixl/gpEvW1
rmxtGpJ/m3Pn8PVCOISQHIdhjTR6rgir4wWlUJQ/wd87Lkbq5T+1K4Gbi/Ui6YrP
440ET6WU6rfeCq4NMvwVtqZ4UmcaVUMJi9bUVhrbZ3omm498tVDzpG2aB8XukI81
fKsHHCnIwqu7sCKnrFMNE5bvhIdryZNdPuL7maMolsfU7qqx5sPHBusE7Za23kQv
XSzQGp9ieOGWUj/ahjlBtbY7KbzRplOJWRyPwVb0X8oAiXkXpqFXz1+YwQZFk/oi
o1dC9RMqqq9fBGWStRFQs9V0pzTkpf3Be/Pluw6NjqQd1InRWTKJqHhIXMnZAwv9
fNckPqv1zq6ONmMWZBCZX9pJe92sfSjZJYcmqj98/fyKIiOa9ze79h3kgjLiKawF
BqL7H0OiVEqaN9FRKXCRkGklCH4D7OfTGn9r5lQso/xZHbgZUg+PPUQy/RCx8dhY
LQsUT9j2KbriqErBFbaK+GdF09aoXz/bm0ndVrmK8/w7vVmBrYUD4yi29n82hh1o
qNqkDjbWARAYm2zJS7ZM8xHitOKK+dlG2uAn57yI4hON6pEHvmQe0/qEKp387Evm
x2I1eV50VtURDEZxFtwCq4Z82yvhv3bq5PNV0wdxnQrG/rx7YKaO/mIaxzyQGAwE
TKTmQvllQIbcT1ve66l1wSck8K/dKlOIzTRBi4uPyJSmXpDqDIzEmp0kioJ647bi
r0SX36tm60VT0Cwb83u1PAwnPArcUV0guJ530Wo5dAAQDhz993OTuDvznhjp5PDl
rlzWFHWp+CGC4Vce17pI3AK8Cjbcmif6qPWDyLBrXRIsOkMKoQs8KQOmDe9Kay0E
u1L3LDFrPvqot/p1FONJ4rbHLCg+iIYpKCzP/EpzTJ5Kk1jpWdolIptsSxZisGJY
3UN+L/wYqNcRQQfcQxzDGsN1YJ/MyYGxOx1DR1LYFQNmEpoY3+NCbySwJbMYpWLf
GeiovoPCBp3tPIlb18gcDVAmAxhnGzhMAnQCuNPpxHQiq/Ql9U7OyO9rZnWiQFoM
isPLEGVk9R+btq4Jou5F4AQ5ePulxs0KMecRMD9ynG0CQ/Tlj/8tmNGVIXDii6+L
BxQEFHPX6tQ3jkDUwpatl9C0zTvg5TTKOTC28wGFAF6WUUAGgc2eLzaCXd0DDnXs
gkX2IfX9FNHDK8Ssn7xBYW/ypDRd92c3iNCZ6VBJRNCw5tQXe3lfrE5+gqjDOhjz
33qKIUTTyK47WkGrXfvnHAflmjEtxg+8P8CW6QiGX+hEjrIcnXx9xb0Qp194b8F4
9f8wwmpjGmG1gPOWfUHAQOYav0XV1wr3FX+6lXskHZnapWerFe5vvYjS0WYkYdju
6+GOiz1naXMdfNmDfTUaDj3VxGm3fMrt2wn3WqjJNIRB9hRXJ3a0WZ9B8CvCmUy4
oEPP5xW1slueaH5v5uFsVoq20KxbXiQWY2taUw+zfaSxFw9DhcTbPrXn10AFKPPi
+bF9yRAyonjqAJ1e6fdHElgSlsi5NtK6dRT/lGyEvBIKvQAr+TtK8DIeR6Zgm/hq
OI1iWvXXaDE+9lHiCeTV8j5NwD6qXc412G7UmX9+UpRKFyjIlh/KVLiWy3BDOTrf
ZR9J8K1rQ0BVNfoCfKs0dlRWiO5P3IKCWYA/P+NxOp/2ckgCxxLSxw23Qe+wxVzH
wottdM+KAHGOQzbnnrN60IdNH/8mroRaoLQpHt3bhRsAK1DIs4zcgF3BY+7i+i0C
VR1TADeKE3xwLaG/Yw4k7bSBFFxOk/v5MVuVwHdLLiqN9rs3LnLpMqnf7hBq5bkB
rJiKs3eYCAtuvM8mZfo1UDk6Pxl6qyVTTAY0L4a08J0v5lVIRRdyUSh8DsVxha6F
awkS630+ZvDxc8j4u+moD/59n8UvTDOKeByuUmUDQd2dbNXr4t4XM+K88pAXK2yG
li/LrrkhiUSfprYS7iNO66PYcG7+cEpq7sACb77MDNM5DPIP+YrMd83iYZ4WxeWp
H+tP/Cg7PFJwUvOy0dr0RU0F8Z7Ii2aisOkJ/L0iGNloltGXTpAOBs8LjggM1RVM
kwg8tdDEv9bwq9ISSE+iDtCkOivR4dv1ZZaNvJeLmhJCpfkXuJUTfK+CSC1kfv1G
CzTP1VZ/zV77kWxWhBDKcLQNLM8EvcY6R2M1/YJFoEWDdZYek3UpxdRn2LYacDlF
juKiXN8DeuA/p1rmIMljDCdMX5Zok2jeVBBg3GiZV4fL/Sag45SIIAh7OzOCP1Jx
F/vHp81upi3kGu33TEEgKXb9aeE2pLSk0+jQ4L3VLIklqSBswauLzz5r67Qhxy/G
aFD5XUtejgsaZoT9Fk3Jxy/0bPmpK9pPuDIFxtfgCNf8sPcTLRFLbgNiaMdgjXFC
84C1qKbOPBUAlcrWY+kxCowyViMOc1gZoZ6YYkPuuiU7OkgOs4sLO+/ZffKDrnOt
FAbKU9YczpOruiHtU1YtzT5/nnWlXUvnt8Kf3+NheL1LfBL9YCPELqxHzr03W1I/
cxIWn8u8WX7IfX7CKhBDEeasdU99tTxMUV/wtqXM7SMccCEt4SQkNSZfsE9N9Dnb
CK/8Kh2p/7tuNOV3V19dLuOTxmbxlJ3QnUtxsGYxTztHeL6xARnnHhDlSJIlQxRN
2bsFr67S367zlSwabZzH2oAsw026DaAdRwd7rP8xoRmb/WslaMJBqseuQ/VZUxE9
NwblGiCePHHtZznMWwzUy8DRVQ/cYTlmPQtCEI+2txj4SsapxPxTadNE+B8SwbD2
D6OH7lTMZ9u6+wglWiu5sqaDWO8qXN2tWdS2s3l1QU4hawpZFQ+6YrKCyNG15Dyl
XM0Xe5AmHyYu3DQg00KBL8NJATtf/ruvyNkjD94hErtLWCKQ/UpVc1B6zS1qN/Zt
IhlRDqhAk4P2Y1bOV0H7Guz7JY7EpqdTUMZIpI8rSZ5njvX0zEdMfIcirXlliD3K
/Pzg99uoO/vPGGj15Z422W28/tvg0MTztBMaf6y39BwuN7cAPHlWgQ589MJFSUm+
hDNmCzsfsK04Q9/JUo8LzBcC4wdbsOGgW0HwichwMsJKVDwBAJ46fl8fxC0BAizB
y8e0QnXWAxgcx+B73Ns4yBlTZAQrZ7AshWbpo9lQsoU6cE2OxcNq94aQQqMXWWKs
8TKPLPkJHF7VSTrbRKcnvOSvHs0+jHQeIgyZaQPJo4r40ozzTjLW0UqSVbejUjaP
t+AEOPrs7T4JYbv9X3Ffm4oN7fzvyr0pGsAX4smqtT5m9bDQoJhoW03jPsryUjJS
oANDavi6xbG04LYlKdSFSb/ErtOBmZPHv6eo+N5hy3bio4g9Zra6Ksi+jiGXJTOz
qiMA6t5uyhHqlNSDsfzyhHnlA1BZvIp8o3WfxOqQQsBmREu8cIPUG5iRnZ1Fd4uH
PLuRgphI8jGEtt2PQ+w7eSNhnXHx4HU1MOSthDUI7wQus0husuMvnySLwUV2O7E3
WuLHzCQ7TX7EmJdKYW6pZZlBwvz14uWLnRVSLRHi9FepFwA/WfXxyPdY6r9EX8uK
2n12a+leMtIG5rHN54rEDB/ThFpawYUd2+pwspkJkDukQA47WPkw4yKbKZzY2xki
PLeo0uMRb+9jBI2WMi6JlCfKapJeKvE462/Ksc6yi+FJgfr5SIvkOoYInaTnIuVn
rwayzMTja3rvIAoOmU05bKromBZBkQrHI+FSNrmTUO01pyT/jjfdWL9F6H/jVESg
EdQ261tL5Ary/mFX4xZgqUUfhKPwP0EbIT+iAb4ZVSsBAEHUIvdM3PrURy/Z08Cp
Yc6Zw07snUHAudEOw1tKxxGztonJK8iXC44Y7EjgfFLpXGLptdvdr6mqBbo8BHFr
XrmxTKd7SNUCfglz4LcoRnSq8i3CNdlSoSyoaU9bYp6OC68eyiWh2YKYcsx1Rp3g
6A0MyFA9wSMe0P7BAeskrUMIle+V+1Gf5jwlr2dd4jj6xB1Qe9VI7wzymVNjNCTZ
8m31cc02aiGIanMF09dn4MrhPpjGpRSW0QBUaRIsDR/JEujrYBaOv/MvovtWevvb
Bx3oPNth9puxX1OELFhXceknyBp3AZ9sRNCkC/IXY0RjzMuHMEbqzCc+ov5FI0UR
ITW2tDI03AcINS/wwBVD61aHVKjDyRhP+ViuUvx0xIbedQi4NGrCFQNbPdvvJeFg
oWOAoI2Xx7azOKZx8DFvjCfGZcplTASCRmnbj6mfj/LDjH/1v+b+bww2Ym7qjsad
jHphTpReSnQHpgs59xax1Qwc94KCDO4BoywkxT6l/tq1U1Jsy5ATYued7ELkiN06
3/lQ/nrqAgvOpwBwHmun9QTSarcYwD0l5MOMFm0MkaHk8pHUWQGOcJMYELdKuLUU
XJ8bWYO31Mvyf/fv/AqHbzBBNsMLlh32w2wW/4vOxc0OqD6x7qTc5G+RfUk2fpb1
ODMJPDhmjbBRqQRZQFg9faBm/gTS9DuBvazvGIhUkSfRc2C9XujlUvMpyYePZM9n
6KmsAMOYugIVqgszYe1Pd7kUrB+dxWtTefE1IQNtjAbVJ7+DaetJh2KqriTCX1S2
nirgbSqPevPGuFJK5uXyeRRfiBu2cT8Bm0NW/9uIKVNaOyzqq6uMTSm1ax405/Yh
XCfKwZ7NvjyoWuAAGfXt5m1C70oCGcvrCF0KBGnGGSvasdDhhh+qhfWeribjXjPO
U0d01J3JIkkqZU4iFzh4es1oKiRP3OgK1PQLb+CSePgV0fgxADk/lzz/9H8Z4p9h
yCh1aGJrC0Vh0vJ2MLU8LICumUzGaMLMp1Dvd8yCeUA54XqjiMHxcmws2pCeghFN
GS+dGbQ2zwjHdogYt4sRgq9iOslT91hRV10wtJ0EmKS+zMUrrS4uyVg9CdOxi4c9
2ezI/BWP5L/AQyuEmhA0yORwGZXwuZhqajk3r48mvYgcC8ZhdiRbsc6GDX+SFW/q
xxpq6ZWJ8VmfS1v2oGR9QGJoJdlphzotjD1yeZvIyite7GE/xGNyd8we5tnIiFgY
CWVOHKAb+0y7iGn+HThUuN9VL8XrTtkhobPYiEu3HIyzRlQTxCC28eslfBkT/zq2
BtKkBUdHzSqOQ8GS9x2zobIYFcFR6sgc9Y2OKvYz6Cucww1qUd6O7D/5PGXIahYi
eYdagh0NQ39NS5NHlA45wAjDVJUkfYdP11vwJ4B3+Njd4ZvRqYfD526GwNK/Okmk
geB+icvLBPlApClft6vMRcajuxf0rLX0Y2VF4B/DAZAqH9bs+dLdsxZaSbxMU+aj
/2roOw/3ZFwRmtsRZCO3q4+Se+10mkuBfS/NpDFX9NQ8jS1aHL9/gs3xCdb+xKAt
WZFsW12IsqqlJDnBcpNEJD59N0Vaoz73m9v4XQdhSGwKbhedz4aYTBgTdNL+OgIx
QZ8+1vnkJDW0SQ1OqACE6/dVXUy9gyLhk7lCnPA9R64lkDZ8R3dh5qtgWXyn/VKI
4rxYOZJJ7K95qrpLZyx3U0inCs6LSb7KFIlgr79BNkGDsfGQYLKtkyhWG9Nu/7AI
X6krAPaViPron6HF1al3qMQN/aMgz31aT/I49P4qrHi5bL5+/iPANF/451WV9+Zj
w4/rfehUCOiQoF7vx/eJzjtrRcHfnwOzl9erNq/b5PJTbc96OVHO6rg11qnxcg0v
yhZoLFNaQ0jcB+ZjW/tNANM5gotn5+8/vWns8IdEEQtmoM59izTJiZI/F8WeqrQF
ksO+hq595RDtgFNSbc0Zvg3A9s+DZWYcozdpRxoAgwbWWQ5/pmjxqK4BkxsMyCHx
WNdJUH5Ho5j/R6v5nXH/Ch8ZGITywtudkgE5hBFQ6HDhkhn2Pf9A1WMaEs+k+yLQ
mU0GyC7ljnUHeXN/DajjqXBhrko85fz5XRyiILVL1VqrA6UeeITGAzAmdYz+fJTi
oEuElo+NvEspwWSEFfZPC3Gmox63GRgW9fRGfzIveu/hX3xhw8NCuI6IiDw/LYz2
1nr7aLuweLHxLDzLQ8rqJ+wNOoOwK7fMj+qXcB8/3be+jdkCmZPvnrdhDDMysNS3
YPt9ZTJRKpHA4nTaP89sSLaQFFI+CPv3JwzmoU0mNsL/9mBtm3mL1mQzuvvyhJP8
vuBfzOyU+U1tEELqtmFOAuybf/EPVIKGllMdURodsURai1tlwomHO6hM/zBuUctC
GWCr04vTObN/eN/O0GZwwx5xEtWWLxaV8pSbCOp5O4II5mygBgkh/JgdgpBlrE/Z
ylO/O7tioqKNji/loyMZECFcviXPB+dsfc/8QJHsxebrmbQF2Vh9r84DrxmNXi7Z
Zag3oXtTF/mqiifNSuNijlsuELAT3spDtkXMKH8tn28mIWwmgm5nnq63xnA4+t6+
5uNls/N2vu27ungBtQ61tIjDwxLtvazaaZA6HXV+mLE26y7dQdXLodQfpHZ3jG4U
kOvxoTer8+/X4mBDiGINl8JpenNSuubiPkTQ/HPHKWDKTRx1u9RrW0wCpHjnJA89
Toy6tP+oTDpkeEI016pUFda5mLBFE5B6NRZJIwE25EiA6ZS8cKvzblAJ/1tZlqJG
NgY/eM+lxjhLK7mM1VjHmW5yyBVK03mvbS2S9K3+jPr8j4Av6qhU4Ojwpd/QQFo5
pEqdBGM8J+WlvF1c4+dNRR6JUPAH99TAOn+1jnGbvKioXvH2sD/4JbfgFpC4b6el
6BhbUlK5eD+ha9tS4eieAQWcg+xdkNmsTugPnxCZrq9jjqVjahV+s/FMx4KMXbnW
u+tyY0eFPF4SI8ulGLhMXKhrkU2bkdRHxcS5T0N1x1cBmB+FcptdqjjtneN3hVAg
dhbmPg0zNbWij3g7CcQF3bpSTLzB4Osg3lphgYSEvUsUn5V5/qpsxzO71d242yG0
pMwIF4zKUqTn9MGeNZvS15kTeUAIejhEgyKaeXXl64lpCNlU1CjugfpA57S/4d+z
JL2PWklWhKB2pxpxX7kqIHY9Jb67DwptvKnU/9Ek6odktx33EGJPiUy4PDIGQbWP
AJKHDhvAO+oDcHLzuEr7HyCzF3rBrYbMhShzyuWEmeUtpysWJcXHX8oToB3OSsie
Oww86nOQoVS4cdLElWxKNLpULX3ixN2yfJWob1h9fqoSuK6g3xv10XaTFm2iUYHU
VmK/galyb3WABsFoUWSLDUs6nK7q+6BI0G5PPWpER8Pi2g557vjC6sB6l8ILike+
rGI68+NqgMduOi4I0vOq47dBy/EvTPVZ6jBum8c7b4Uxt4vdcX5wTPfmv2ntSmH5
bX1VmjnJMKNEwSc2ul7Ygubta4L1oSh12EuVsqvOYzS+uyR8XaUbOVh2EuAZa7Nt
0BLxVDAnAzzNKBAW/XlB70WAXHqXdOYinuae5bXQk83OAmviYmh4ktlSnkXi8Q5n
gjwHWlUV8oas6bsYI4HXhPrF2OENhINGYr9+e4Q24wnzh2dN67s5jHv/EyWUMZxf
R9X6TYJb4e18+yJyFoRDXcxLdPQfUH6Ebox9hWKDUrGQmcskC83Q4r9XXijdCWp9
P9zUC71YLwFx5fxYL4k9gFWPZdpyiGB290bHt2ENBdGtDAQXm88b15jDKoCyriMB
wdpimWZDf8LGRm27My+aIeSbVfJbu7Sp4ZtT/n5ssj/wgp5HuIhacmW1x0jCmJJx
ptGmr2xqhLyYsyUIqjpH/+dXtWltomMUrevBJcSHw58oKFut0pp3GHvdpIY16aWQ
NQc1VSbX3xzJWt0vjEYxuGk6F8Uu9PAPDheHO4UrpJ8YzClfa4ZzEa5sVj3y2P10
ueT163YEcum/x85JbVaJIatzetsVjji79xAs2wbWakxmF8ZJwnUAjQIcC7gCFDYp
4o4l3ot7sgTVJ4ukmFqOSEDS3rOhrvx0F+zb6rQi1bXho6P5aWWPnIOiEzVoA6hd
5Xmk9NTSKnTiNYcrNzn8MK/Ho4CmvSgveZpfTJC9ZIteRKVjPR4q7d55vwKvO28h
gOPQrazbD64cNYDfuoK+h53FrpUzuwFHVX1dgkTQ/xxJKuWTmAfv1aLBI02Y5tdF
gEXR8R/pF4Z9xbG9fiSEfTzK60+yrtpFYExnrJxA7r6/87CXvM9wdW0wRUkpfjA/
R8NMuf7h5buXVF8pJS0UEoCkoS8sLEolTBUKlx/88HD91zOk3+ngWGD1djejdVkX
Vq8/U3uTHk/5EJWVQlkWS6LO6uRAfBWoJ/o+SGK4yrBcQrF/MgRuTagE8VJYL0tz
9An8Mu89l2EJNZydR5VkVqRSkoLA1wS6RCypWVDmobjGFOixF5GWqEP0KQ38A60e
axgA1INQOUKzVwjz/paNCbJz+aoF8iGAxuOlgjPStkCtA+B94drGlEXdJRR4iX93
/ZkTcmFnXdTDjW9beo0i9RbdX1mOhBMLYJ1c7gLs/sLEjymrz/iHX/XoZguFZ8w5
VhJGMsf657WP2SqM0bcuCNqwsCH2pH+MheY+tX4P8btCku3/lAkKqXcGn8ltLaVA
TFzuD5CWLKiGQp8kP6cPFstrMBJCKXSvfe8jaTBvGAWWVvVXoTycqt+mOAR3Efb+
KrY2q5DxjlBh0HNzYareeNelKhgTfijrDqfabkxW0IaOiwQl/4l4xHh41R/xo6pB
dFE8Az26Y9JrIGRQ9yZz4Xxja92b7MA76fPVXOigjLlqcpI5SIw9kB63gE5jZBXP
nnjKX/OxIjpRXTvl252j2lhj0gnD1radcErBq2Vg3DC06Jp0ZiiabTILMrkbWUfi
zD829/bVr4shffKfp3f6quMgdeZBoHYmqMZ1EHF1HG2FGxx5D0Ptd91YBrEj9blP
sqCvnTMFHJFZBfh2jRiDMFwwBaiEI0OFdz1pv4gQ1geSoAFUyLofjZ0xRlClbnVh
78RCpuj71D1ESPy/XHq4x7wNyZVy7jofn5OhXnOTfNc=
`pragma protect end_protected
