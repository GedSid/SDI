-- megafunction wizard: %SDI II v15.0%
-- GENERATION: XML
-- sdi_ip_ii_tx.vhd

-- Generated using ACDS version 15.0 145

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sdi_ip_ii_tx is
	port (
		tx_rst             : in  std_logic                      := '0';             --             tx_rst.reset
		tx_enable_crc      : in  std_logic                      := '0';             --      tx_enable_crc.export
		tx_enable_ln       : in  std_logic                      := '0';             --       tx_enable_ln.export
		tx_ln              : in  std_logic_vector(10 downto 0)  := (others => '0'); --              tx_ln.export
		tx_datain          : in  std_logic_vector(19 downto 0)  := (others => '0'); --          tx_datain.export
		tx_datain_valid    : in  std_logic                      := '0';             --    tx_datain_valid.export
		tx_trs             : in  std_logic                      := '0';             --             tx_trs.export
		tx_dataout_valid   : out std_logic;                                         --   tx_dataout_valid.export
		tx_pclk            : in  std_logic                      := '0';             --            tx_pclk.clk
		tx_coreclk         : in  std_logic                      := '0';             --         tx_coreclk.clk
		xcvr_refclk        : in  std_logic                      := '0';             --        xcvr_refclk.clk
		sdi_tx             : out std_logic;                                         --             sdi_tx.export
		tx_pll_locked      : out std_logic;                                         --      tx_pll_locked.export
		tx_clkout          : out std_logic;                                         --          tx_clkout.clk
		reconfig_to_xcvr   : in  std_logic_vector(139 downto 0) := (others => '0'); --   reconfig_to_xcvr.reconfig_to_xcvr
		reconfig_from_xcvr : out std_logic_vector(91 downto 0)                      -- reconfig_from_xcvr.reconfig_from_xcvr
	);
end entity sdi_ip_ii_tx;

architecture rtl of sdi_ip_ii_tx is
	component sdi_ip_ii_tx_0002 is
		generic (
			FAMILY               : string  := "STRATIX V";
			VIDEO_STANDARD       : string  := "hd";
			SD_BIT_WIDTH         : integer := 10;
			DIRECTION            : string  := "du";
			TRANSCEIVER_PROTOCOL : string  := "xcvr_proto";
			HD_FREQ              : string  := "148.5";
			XCVR_TX_PLL_SEL      : integer := 0;
			RX_INC_ERR_TOLERANCE : integer := 0;
			RX_CRC_ERROR_OUTPUT  : integer := 0;
			RX_EN_VPID_EXTRACT   : integer := 0;
			RX_EN_A2B_CONV       : integer := 0;
			RX_EN_B2A_CONV       : integer := 0;
			TX_EN_VPID_INSERT    : integer := 0;
			IS_RTL_SIM           : integer := 0
		);
		port (
			tx_rst             : in  std_logic                      := 'X';             -- reset
			tx_enable_crc      : in  std_logic                      := 'X';             -- export
			tx_enable_ln       : in  std_logic                      := 'X';             -- export
			tx_ln              : in  std_logic_vector(10 downto 0)  := (others => 'X'); -- export
			tx_datain          : in  std_logic_vector(19 downto 0)  := (others => 'X'); -- export
			tx_datain_valid    : in  std_logic                      := 'X';             -- export
			tx_trs             : in  std_logic                      := 'X';             -- export
			tx_dataout_valid   : out std_logic;                                         -- export
			tx_pclk            : in  std_logic                      := 'X';             -- clk
			tx_coreclk         : in  std_logic                      := 'X';             -- clk
			xcvr_refclk        : in  std_logic                      := 'X';             -- clk
			sdi_tx             : out std_logic;                                         -- export
			tx_pll_locked      : out std_logic;                                         -- export
			tx_clkout          : out std_logic;                                         -- clk
			reconfig_to_xcvr   : in  std_logic_vector(139 downto 0) := (others => 'X'); -- reconfig_to_xcvr
			reconfig_from_xcvr : out std_logic_vector(91 downto 0)                      -- reconfig_from_xcvr
		);
	end component sdi_ip_ii_tx_0002;

begin

	sdi_ip_ii_tx_inst : component sdi_ip_ii_tx_0002
		generic map (
			FAMILY               => "Cyclone V",
			VIDEO_STANDARD       => "hd",
			SD_BIT_WIDTH         => 10,
			DIRECTION            => "tx",
			TRANSCEIVER_PROTOCOL => "xcvr_proto",
			HD_FREQ              => "148.5",
			XCVR_TX_PLL_SEL      => 0,
			RX_INC_ERR_TOLERANCE => 0,
			RX_CRC_ERROR_OUTPUT  => 0,
			RX_EN_VPID_EXTRACT   => 0,
			RX_EN_A2B_CONV       => 0,
			RX_EN_B2A_CONV       => 0,
			TX_EN_VPID_INSERT    => 0,
			IS_RTL_SIM           => 0
		)
		port map (
			tx_rst             => tx_rst,             --             tx_rst.reset
			tx_enable_crc      => tx_enable_crc,      --      tx_enable_crc.export
			tx_enable_ln       => tx_enable_ln,       --       tx_enable_ln.export
			tx_ln              => tx_ln,              --              tx_ln.export
			tx_datain          => tx_datain,          --          tx_datain.export
			tx_datain_valid    => tx_datain_valid,    --    tx_datain_valid.export
			tx_trs             => tx_trs,             --             tx_trs.export
			tx_dataout_valid   => tx_dataout_valid,   --   tx_dataout_valid.export
			tx_pclk            => tx_pclk,            --            tx_pclk.clk
			tx_coreclk         => tx_coreclk,         --         tx_coreclk.clk
			xcvr_refclk        => xcvr_refclk,        --        xcvr_refclk.clk
			sdi_tx             => sdi_tx,             --             sdi_tx.export
			tx_pll_locked      => tx_pll_locked,      --      tx_pll_locked.export
			tx_clkout          => tx_clkout,          --          tx_clkout.clk
			reconfig_to_xcvr   => reconfig_to_xcvr,   --   reconfig_to_xcvr.reconfig_to_xcvr
			reconfig_from_xcvr => reconfig_from_xcvr  -- reconfig_from_xcvr.reconfig_from_xcvr
		);

end architecture rtl; -- of sdi_ip_ii_tx
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2023 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="sdi_ii" version="15.0" >
-- Retrieval info: 	<generic name="FAMILY" value="Cyclone V" />
-- Retrieval info: 	<generic name="DEVICE" value="Unknown" />
-- Retrieval info: 	<generic name="VIDEO_STANDARD" value="hd" />
-- Retrieval info: 	<generic name="SD_BIT_WIDTH" value="10" />
-- Retrieval info: 	<generic name="DIRECTION" value="tx" />
-- Retrieval info: 	<generic name="TRANSCEIVER_PROTOCOL" value="xcvr_proto" />
-- Retrieval info: 	<generic name="HD_FREQ" value="148.5" />
-- Retrieval info: 	<generic name="XCVR_TXPLL_TYPE" value="CMU" />
-- Retrieval info: 	<generic name="XCVR_ATXPLL_DATA_RATE" value="11880" />
-- Retrieval info: 	<generic name="XCVR_TX_PLL_SEL" value="0" />
-- Retrieval info: 	<generic name="RX_INC_ERR_TOLERANCE" value="0" />
-- Retrieval info: 	<generic name="RX_CRC_ERROR_OUTPUT" value="0" />
-- Retrieval info: 	<generic name="RX_EN_VPID_EXTRACT" value="0" />
-- Retrieval info: 	<generic name="RX_EN_A2B_CONV" value="0" />
-- Retrieval info: 	<generic name="RX_EN_B2A_CONV" value="0" />
-- Retrieval info: 	<generic name="TX_HD_2X_OVERSAMPLING" value="0" />
-- Retrieval info: 	<generic name="TX_EN_VPID_INSERT" value="0" />
-- Retrieval info: 	<generic name="ED_TXPLL_TYPE" value="CMU" />
-- Retrieval info: 	<generic name="ED_TXPLL_SWITCH" value="0" />
-- Retrieval info: 	<generic name="TEST_LN_OUTPUT" value="1" />
-- Retrieval info: 	<generic name="TEST_SYNC_OUTPUT" value="0" />
-- Retrieval info: 	<generic name="TEST_RECONFIG_SEQ" value="3GA" />
-- Retrieval info: 	<generic name="TEST_DISTURB_SERIAL" value="0" />
-- Retrieval info: 	<generic name="TEST_DATA_COMPARE" value="0" />
-- Retrieval info: 	<generic name="TEST_DL_SYNC" value="0" />
-- Retrieval info: 	<generic name="TEST_TRS_LOCKED" value="0" />
-- Retrieval info: 	<generic name="TEST_FRAME_LOCKED" value="0" />
-- Retrieval info: 	<generic name="TEST_VPID_OVERWRITE" value="1" />
-- Retrieval info: 	<generic name="TEST_MULTI_RECON" value="0" />
-- Retrieval info: 	<generic name="TEST_SERIAL_DELAY" value="0" />
-- Retrieval info: 	<generic name="IS_RTL_SIM" value="0" />
-- Retrieval info: 	<generic name="TEST_RESET_SEQ" value="0" />
-- Retrieval info: 	<generic name="TEST_RESET_RECON" value="0" />
-- Retrieval info: 	<generic name="TEST_RST_PRE_OW" value="0" />
-- Retrieval info: 	<generic name="TEST_RXSAMPLE_CHK" value="0" />
-- Retrieval info: 	<generic name="TEST_GEN_ANC" value="0" />
-- Retrieval info: 	<generic name="TEST_GEN_VPID" value="0" />
-- Retrieval info: 	<generic name="TEST_VPID_PKT_COUNT" value="1" />
-- Retrieval info: 	<generic name="TEST_ERR_VPID" value="0" />
-- Retrieval info: 	<generic name="AUTO_DEVICE_SPEEDGRADE" value="Unknown" />
-- Retrieval info: </instance>
-- IPFS_FILES : sdi_ip_ii_tx.vho
-- RELATED_FILES: sdi_ip_ii_tx.vhd, sdi_ip_ii_tx_0002.v, sdi_ii_phy_adapter.v, altera_xcvr_functions.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, av_xcvr_h.sv, av_xcvr_avmm_csr.sv, av_tx_pma_ch.sv, av_tx_pma.sv, av_rx_pma.sv, av_pma.sv, av_pcs_ch.sv, av_pcs.sv, av_xcvr_avmm.sv, av_xcvr_native.sv, av_xcvr_plls.sv, av_xcvr_data_adapter.sv, av_reconfig_bundle_to_basic.sv, av_reconfig_bundle_to_xcvr.sv, av_hssi_8g_rx_pcs_rbc.sv, av_hssi_8g_tx_pcs_rbc.sv, av_hssi_common_pcs_pma_interface_rbc.sv, av_hssi_common_pld_pcs_interface_rbc.sv, av_hssi_pipe_gen1_2_rbc.sv, av_hssi_rx_pcs_pma_interface_rbc.sv, av_hssi_rx_pld_pcs_interface_rbc.sv, av_hssi_tx_pcs_pma_interface_rbc.sv, av_hssi_tx_pld_pcs_interface_rbc.sv, alt_reset_ctrl_lego.sv, alt_reset_ctrl_tgx_cdrauto.sv, alt_xcvr_resync.sv, alt_xcvr_csr_common_h.sv, alt_xcvr_csr_common.sv, alt_xcvr_csr_pcs8g_h.sv, alt_xcvr_csr_pcs8g.sv, alt_xcvr_csr_selector.sv, alt_xcvr_mgmt2dec.sv, altera_wait_generate.v, altera_xcvr_native_av_functions_h.sv, altera_xcvr_native_av.sv, altera_xcvr_data_adapter_av.sv, altera_xcvr_reset_control.sv, alt_xcvr_reset_counter.sv, sdi_ii_tx_protocol.v, sdi_ii_hd_crc.v, sdi_ii_hd_insert_ln.v, sdi_ii_scrambler.v, sdi_ii_transmit.v, sdi_ii_vpid_insert.v, sdi_ii_trsmatch.v, sdi_ii_sd_bits_conv.v, sdi_ii_sync_bit_ins.v, sdi_ii_tx_phy_mgmt.v, sdi_ii_tx_sample.v, sdi_ii_tx_xcvr_interface.v, sdi_ii_tx_ce_gen.v, altera_reset_controller.v, altera_reset_synchronizer.v
