// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:11 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qjKBZe1dy/dA2iYAJr6Uu+w7kBTUdrDpGjVDV8XYq2CQXxP1bqBVi5dQt0Waadpb
DTSSMByYI1WPR6DAz5PZ2MdPQuPm+t0EeyS6Vo+ieUjDZY6n7QGqNeLl7ENnfP8G
tuQbSTb4fESjxtbPRfGnW0pHVHgA1O4g6G/EOXF6iqI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15968)
V4kOZVH5jc5NjccjCk0NM/jaOMUMxajOYgAaCUQPw4Ct9sx84rocxIpj1QGIDvCL
OwogSFwZLEZAD7tFbHimdXC2SmU0IdMRW81sWD1s1wAjz1tInQy4+fYbAbyEQ6EC
dwl9XnpV5HY8Ep40kAHGoE/AChduhNwOCvj1DO5/ueznQCZGMwVV0zeNygycDW/i
F34Qw4Db7iQo7o6uoDvkmQHityfmNiak9ApLB6fHE3CrpgV2LRFdTarnvi5WXrhj
YeUGK4+PLUyinjAU0unqFKuctLd4rgYXEu6byNL0aN8tRFc0k9Ga3iMaDt4ka6d+
0OHED7LTtha1Njclll97eoT7iXud261DPAPXahVgnZzwxeFWpQpbCStqdukcr7Nk
wowFsvJQqDSNsjVhvRkVZRFCvp69yHY6gQzw8VmmmHdc5k4cNyPhuI+rUP+TK2ta
33vkuw3aBBO0H8Be5Gt1xXaBalJT35blaDRmHbIHanzJkqNHPy310jeszt98Wr5S
Sj2bAJ7GQWRPmu2BTiItXP76i18DbRj0rJ68PGtaTWPKXhX0yg1Pa1xXC5iuurnT
CThzHojNxzcr8NAlTav/7KJFxSDBS9qznzjvtysdrJ2cLXnnGnrpAi3RBFtua3f3
KWEc+wYTl/UQIsEZNmDsm8d14CFXtT6m4RMmuj/EVfXqAHo5RayomIrzO7fqo64M
xK31zfd+KIYdCBoJOyD43GQtRGWQYYXh6QFhHdrghvO7efJoubcyRFl0WnBbeYA9
emD70f+omXoFlfgemzVBWPs2jHRKwxo6imDp1lZVXFjn/q3Bte6YZnr0nWgTIlXs
O580aLIIs1LLO1jv2ND0AfcmmXnHuEDlH/RlQjbF1ZUsLyzqxYErkRbyZikGMHd6
ELGqKMI9DWj39xQyc7ZHQ99ZeikTRTWeL/WbJzM3EJlE0dBlTxaGF4WD0PKXQFY1
lo009A4JRS7252epmUxCqLBpBiEYIvYJ/nufc7x19ZONjJYYWWYAYmTh91gkwNp3
vwiIh+t/taMltBFGfheIh3ocsRe/0Ai95FJ3Tcq6mQoK545xO+Mw74DnfyDPlO4+
kEaTi1WBvy5wuzMkqhdfdSaLnnxZYN7hj14JG3lb/sM5t/tSa+Iafq48+cO0Nix6
Gteyp6Rw1xxGUxzUXUEIWPyEEYXSZJ+grBIrDhuFH4yxVjbgSs2f+CsaAanBV6uQ
lZM/XGRY06S/jpMfxyTuRNxnO1GbEanFM2aEiPA5JclsIeZg/Xl++OytaN5j8S4w
/51zRgzobv35zh5sbVqPvM+UtGVRBypuudc/eQFKrZPI02z8S5a8Otf/Lv3EA56a
ajbzYEChPpoZ2jsZx6BY88q0D/dRrvMroHqUKq4tX8PGcqhiLODngcP2e/zRF3Sh
QZbdJd/HJXvJTW/VUh6fBAzAlZURwEUdguE8tvw0t8xBDb7s+AdEXV6/JjdeFJKL
T2xiNNg6o0fo/U7FFZJElsCT6hYjH+bQbeyt2XwUqGvvAMSk+nTrsmRihMKGxx3A
WIIPVYge8tNABUCOtBSJxo0BVuF21T0ASmlDnQaZgYbLTzSH8l9s0n3Dk4fW2yNQ
9GnnlW0dciiv22Edaff7ftolSa9i3IT+zW0cuJ1DZAmGT7yOa7PU7QF8R6/mEgHu
PoKotRTFdVmRelYS0I79iJ++MOwI6uQMdczPGYV1Hymsgs1nD2VURrMy876CpxqL
VTEQuOFIzMLtt6piXjkMnNgpUeX2CSGhpPwSTEvzPSH/ta7rHApph0ocfdh/6jdn
7AOyhI8b7hHcAEAqhYfrt55mThC/rhAJwEaZ62QpGZhksrUZSu8I45dg17IbzNbr
/bhE8NHVM//DtNUlMV14kNkYK93Jgfsk025GpsFxxyw7iNkmGpFKRgblfG49Abrb
mxJ+HMPua89dhy451zci14nanQzPEp3K89/b13ePNOX6IikgQ9KXZOL6o06sYSkS
+xHQlAOp6Eo+1R/M/yDL87OTSqmucSsW8na5npHGfSfLIZxj/oktcBy5Ise0E1y6
R2TeZVW/mg+oJowWnALl1RmQr4/pINdjaUy/kv0QTN6gFx89PzuIPX13NRZ9sxk2
ejQ1ccJtSQ1ZoMUABCWSrz90jNA4hJP5IzouDIMCo6W4PgaBTcXAFwkhN6ibwEcU
gjOmdOiJmd6JET/SH0inCmOQ4BzE6UoVZL8AzBp04ylfRQNDODJ81C6sb24hdwol
4/KtvDvE9op9qUbUd95L0NHdfiun1dtOebN2CaW2x9DFx0pZszf6szh6FrMBx5s8
bhZUhtsE+spRMGfGF/QuOlkPzG69eH+HcV67pU1lhLsPOVU/ZtGsI3rUMdka11EZ
BA6ZwoqRiC7AfN8WfAmg2L1ZPLDWMvlJWYkemv18q45RgR0uFT4gMtyBUmdZ6Xz7
LBHNwsf5XyL7p7p6rwBvclXVZg3Jpn6WDgUQuHWGEhUsswWov9x6Zd2mgIsXa7gp
LR8XwLfhcQvk8MLrHXUd2VZz5agX9JQLCRcPr1//FoWqxustgUwtmDfzHBpRG4Ry
t9fs8FXDAVZX5DAGKtOJxtgUjj5X21RKX6cyRiSTeyIPEPLoMj47wP35QGZ+AZYQ
0EnIVjoUwFxGbfJTwKv6P3ToqXG22l2PMXsQBUh+hQU1AbCrDdYQ9fym5oJprEna
7By+SJtlFjS+0J/hjFhTC5Ybg2nwj8LgTpRd+s6Suvf2R/D0ttYufWH0SATIZF74
RR0xAXzv58RVI1b1madOcZcPmKiYL60IGTPQRkm+3V7frUae6sNmkLY3Cz1ee8fS
zYn7yK5lLgYnsp3zjrHJk+pFBfLaAvkn2TwZLSK+S0qsAGAcyCOanUDl9WxZJj+O
/f7Y42uCI1yo4b6rMB4xLbNWLP91S37o2Sjn2Doqnh7IFdKjL1US/SAK/Dm1A8x6
djWYBS+LQj5TE1cnvdVbfzs8t5WRt/9ATpVKagGvxI6q7rPbR2G86ZWFqi54DcXZ
8yTAnm/lTkG8rL1SHzudwcrPoQYXYRrE1uTLqUudG+MRpF9pcey5aRfTxUOxynph
nGb8arIqOEXVGrlc8umgB0kdpalZSCFpFTylQJjUJikRCmz1DRKaMQhK7S99yaF1
6YOOt4e5VIz6TWHvoqM+nDg8BRwiVdbLVxYcyyBEiAxhh2IZxwtb/ivE3KoeUVo9
Ahc07f2kX5cZul0ObkxmBMrPyMFfKez/CSElAx0Y3WohdZSaS3T0wyYDjXA4Ap7r
qeLA3k1k0NzP8tqtWUDBs90H7Is/kJ/ZEHLPuVZMvcyMOu+lrYf0ol9mgs/RcxZh
7IbCwKTpHA7dQYiiw4dF3xSZq8o9ksY5gV8HC3bMKRes/c3k0h6M3nsgoVZgTgJW
1bdc+fu+o3x5gOKjuU/sYWlEMqvDwCfPtbejrwmc2WUQx7HOxrVlsn25Sw+rcWmG
vzjLnw8/msv0hJE+r1B820ILKMCzvtHdg3avxvofWbstz0llZ5xgq7kmuyN1qTn6
9m+jW3lEDQCXG7K4tI2vZinmKxek/yQkzVtJD/pwelPsqoAYVDJzlLS2fC9xya8c
L+dV1EWxse1kYPsfPXN7s52RjHHhaCHvuOGO039c9iSxvs/EQllL7sp8L39b9ON+
KTH18OmpNOv5aWB8jxB7TJtAa43ds9zs8LMHbuutpG24/46yubPqfmR6W8KJJ8pO
//76p4Rm3rXpl7QPLT7Q3Mp3vf9A8WhZRYFKyyBCn4GfWc7pD9omPexHY8p5dnO8
0ABsumAcEpHdUCWlhRpkVGfLb9fZRzTYmmy09XNiVLqS6YTIP7szXyFqHHJkU94p
8n/OjoelnPK4A/6L43rV+HFROge+liu7PYxEa+ygbJfZqJ+OHnPOxBwDdoVhkSlL
99RKzXfpD5RrolLI85fdNbjpoTPdAT5Emm7zoOdFRrT/7ccfho3yoH+gq+n0vqmi
TbysJflmBNf9JYplrAZMWjDDOSYqjbotWUojCWBb278q/+VJq8I7uENq/KiaaDiW
JWso57NpLfEWglYyVFrMAle75r2YtIJS9S5IVQ3b22F+C951EAQ9MyDyt4ObBDhK
u/MFwo4/3RGhHP/gJflTpdyKO79g6tVE2JjZnSaRJSpvYP7hzz40XkJbNGXDBHhR
bu//FPh1gBLAcyvzv0NjvFuZNhebzPrcX8vv7Ol7yTx59yuYQtYJkTJNkgcA0NjN
EXx2kiZQctM5/KInURE3BCbhoKeuNf3lrPmel/GQCX7nogOgGNF0VT+35V76xMyk
yyiLW1PDTQt+Pcgd7SlVoGVaOncMSZOLYZkF1J9IyRnPtB5IQTHsKdhiXS6vvb8Y
ohLk7kU+iUiNewPYH/MesAot/XTH3XFVNlUVoUT7U2UFmGUU9YLuTrGlQwBssTKU
u0nowGlfu+YF8maKNjLHkAPhs/oGYN/bHOtmLotKIiKnyKBmqG+3e9zcwRgqcD26
VHri0LenxljoXa2x/sIy1P/YeTqx5NEnOHSmrM6d1HI+5guC/fLuKREV4128GSwJ
pCVBTCeHWpvRl2kooXv0hYUUZkjbjLwSleQLO0o4eEKJLM4HYAr4Gk1Y5+hNxdtO
KsrYpIhIo8IjnxWIfjsyQvZheG1035Mbx7HdM+w9bQTsrrBriwvYZ8hYD6S1Fr2K
OC+356xdTNKiMzTUe44uh73OkMpPmO9P8ocWdwdEnZzbILtRt5Z4C7G75D9OF/Is
vwuU97h6l4gbBbFPsqZ/bERZ7SfiDTg193Hl03fJo+DSMwcyUHD2zfWsRY0HU5cj
R3JmlMBz1rmvxgX8r2TFuQkEXjEBkms07yG1gCR6x8woC339xGzMhkHquu9dKqlZ
+O7iSIn4Q4AmFJ2MnGXcEzrMFKPmT6xOT6ujrjWogCNPNssh6wbPizgOSy/TzwZ2
CY+dgRXqkQJGnSHSwrN239fvdW7+Wk9fODQpRkHVWeN6RwlQJ7Ip+9LjxEevvf2A
PBe36jK9IZ5N763m1Q47t6TTWeHaec3ZP3SqnZkffYBnAIhNpQlyN/hPhGX1ZlTn
/xHGhyCIv6oyLJLi4eWhqhm/gY9TE6jsiS8rS4RTIK42+M+i1wViWs11ACL+HENF
Coh0K5vS5yMEU/6Dg3bFjkP+W9/dO3baC4pz8KGBlhYufAvGU6ny8XJ/RgIj5LiG
Pn4FnUJ++xu6QYsrtP14DLZL1nTiS7dQoi35tzDSSeYJZ5Df29LlUj0VxeCFCe0w
TX8qMv/KyObmnGMFeZ9COVvryXUMF+bhp83Scz2hA1t1+tR56Rkd4kkB1rcSCQYg
RGJXQlP0i0PJOEq7LrQZSDF3DthXDhE6yZCI+eY4lJ8StUEU8RZtJRqAi3ztE3S9
WeXXmEX2ad4WjhQ/qxlz+I4lOzZCrZqi/zVXIimXi8E4LuakcG6mIWXVkFUliG2c
gm65dXHKwrlcfmUTy9t2nIZWrUNAOIFq+qL2KAf6pQZ2FbEMVUrW+cFvXdgRW+I3
JHKvPovlnBvS62neRN8sxz9iXbH/c79sMpX0l4vNE6bC/niAWf8/KEV5kFreZ/Gp
JWdA399mmvryXIUcymCSEXmOiQMDSdLfU1yfYSOQ6Y8NLKdcfTh/xrKmRgb1IBFx
G8qiEYIaS4cGADJ0W11N1GeYWQnj8OJynAMJFVp8zudGlFYi3VvXmXm3DStHfXSW
z2YOWhh/PJfvtxtbN5O4PUGnoKWrKmBUdo+UxKQLgQK0bzXsC6oP5zhB2Oo3TioH
bA/FkyPFVPARyq2M5eFtCiv6kCkMv9H964m/ksdnE51ztdalslS2Wvz5NdvisLmi
P8M8vuY1a4V1dTgBWEwvs25lV+F0UNOmv/rUdreDs/9P08/tgB6opILPp2wab27s
XpIwUhx/piyMKwPfDsckvDUC+OzGKNDOiLZD5oweqHFOPBVxlwGod8nyHYT2P+dP
lYY7GLdHMyI4V4tY0+vFOkt6D2psBQCL/OLejyNJGoNBPnTGtHb75Gpz3jQeqfrc
Fd/oow50ILRs0i0CYSEFr3uoKv4s7CotgdE4SUNpxTr2YShGif7X9K2sD1eYHs5P
50ZxRG6EzQvNYlhYISDH8EF/hFz5PweB1LwjR6dgggv62lOtDhnPaQcc0a4DKq9p
fA2Xz2Vfr4O/QB6FsD/pLffPkGCtnyqrClwYzOlclV/duigCvCQA3Y4QCf4577K9
cNQZPj2Tk+T9r7r4gY/lSfqR6OKdStIcAwFBeTGkjoRZ9D+sorxnXq5G75EeQTi9
lqrrHXDNw2IErny4035R5IkOvJIoEoGc/seG8IGRFf2PdM8NArwvUlwlsPl/EzGf
0zQSqy+CQ5vIZlgXn5+NrM0r0n8bV9zHO2HrH5q6OW0JK8gN6ejUB1AArROhEZF9
jmDOlUPh/2ShhQReLRG5S9fKVrA5iKYW20p5UQZIfCAXaqk8dX8xFCYOSaystcrS
DPNL43hYonDKDY/hg4aht7tOLLX8FxG9y/oaLPGDh5q/xYf1oKIAoHxaIs6g/MJq
mnyUMoNJuwA68LRn7HSqWBhiyqBUv3CzZwYkhv8Ni61ZQkoH7QwAn17y8RVoPbo9
0kP6KRwwNe0wHwbyRFuxe/u18FR5gzt+GlsWbNG7i6btVxMjsEvHetnScOjxkBnX
jMQJt+V/jHtYagB9dOTIj2ixzcs7rgXnnHAIUldm0iTfgdrDwTNT0vwGc/2GCArb
Vas2ubTG8Z+tERBt00cC9qmxgPJD+4fKCeHf3q6maRjWEffxWZMy5N5YQV9m1KTH
AVavi0JZn9G8gWMvZyu+6vL3PdFvRzqURUB6i0OPWVdcg95ODuYKDGJvKjRtWCst
Q+s25UQnJnexwVo1+i42GJO3ylwmqy34RI8UHEBc/Ra81QEubTC7lCsGLruyXWQ3
+zX/OyPIsgvp3Dhj1x72N6uUzHOwxg8futb8abQdbwX41jwVUE8M/agxkyW7b+OF
rWD8cvkH3Xc8yf2abjYzdNP8iEOsiX2s08wNAzcyepookoM5ItZLa1IbZm4lIcMB
GmRH339aFSmdaHQHk//gxK+2tru5cKyCfKwtA8vw04Ys9MeRU+ZBalJ3YJf6gT0v
/RIDw4pOwR3/JlATSIqfjlr85x7082b98D9VSXubhA/BgdS9cdOtQ0Zgt4HXj0dY
qz4DkdlMSjZZmNn85Lji9Dv8TWkTC1vACOw700MRRgZ/5CBQy0GwT+t4uzHWEWcy
Bflfdf6nlAm+Nd/0kIAE31YpNx1hbJmaLyPWjlPfH6TjkgBfcSa6vVuHQsuFv71u
BoT/3geib25n6pBp/NouFYRK7viLBYCZgoaFlNELhjpKgOo7oMxcjIGFDRxkyzSY
MfA4urwkT8J5DBrIqvOCs7Jid9/KkEvkrzDyyolvAEAEl+LyP337eyM7R1E+1dCt
bhcneFZ0qPLvAQbGA1No/QlHo3tjR83lf/GMcfd30ViLGlEKaTPTpcT+ygrh0Ifj
Lk7mXdcT/aBwyK+n0w86Tp5wD0McrlmJeMPA5U0TTROGIiJ8vkXc+VYDlyarLujz
Eslyx+wYcL/0JkGvcIhhbzTCBVOucVtmP1xhiWJE59K7dAmPwKw1/ApY1ZNyeN9c
fVqhIbZU0AzIK1JmesUIF8xIIm74SfROPcUYeonLIYCVsHquBI8OulEoYRnqtl+/
+sYLasJwf+o79SvzVEP3oCyQHQARumMySolTIKV8rr+e7m+wRbzS9jqR6u0n8lYT
EzPBeuHks+lPmyjfyAZ2uzexYWbg/eTQYNU+qGBdkwz5Oine4Gd6yiU6kVmqMLPC
avAckhsJrUTUG6vAQUFynQNkSBn+7fJwjT5bNiDgaLXlGkMvue4aPiFAs211ZM+H
5nECmDMwUo71g3x4I5aXM5u5su8pAvzo4ZQ/3EMhS5S560lmwbPql1B152+VBPrN
LroZvB+NINRmtPyTzkyCDqdt4CfU+BShpL7kjpJRV0p1BWmIMlnHTb7QGMe+Ieix
Mhmn/0HC0Q2s5PTsIoiR55RBfxWFaYPvMOnUj4JoF3vQCMKM7xx8VlerK9yUesVA
jx0q5RpPeiqogzaOTzthUhTh2jPO507cfVJVXF59GOoocZfwD66jim6kNPwU8Isk
f2eTLcDrD4CYJDqfkDBhjUKYQz7vvCcVqollLyZqhPl0xsCcsCPuxGXdcPmkzh6f
BLwHmOciWJvAia0C8FhgowRovz5YFHUKKSqWzKPesU7V7lna2Tewp1YnBBJU4k7o
6DBwvrZzhHqjUNdwrVITgSfKNEAWXgZaJJc5kXNDK131d8shuoX4V/jRr/NlgtGj
KED09FZcbnnuven+j8BKZddRg148nMERi9bGGh1zImNOXjlGJtHUl5Ied0Ddi7XT
ErY4IasnuFLyTY4JZ3WqfdWY45jzv7V8HpTTRqBKyVoC8M7iZJWjF40QE6svwVx/
+PlBbR0hvuVy4Ie8orLGXXi3lFru56zem2u0Dqu/E9KHnQXR+XrhNfj5BM5qxkF4
vXr88qJ/xTO3byudwqr5xQccK5haobni6bf8ucsq+9Ry1mXS1BXasQPbm28yj/ad
VnMbgOBzAlQA5ysKXdfDM8vfHU7iEfsjtCSLzodl1bMchAZ+9EkPpRfhREoHo45I
qE/EgQ1uLCvX6ISulNRrUi3tdWIXai5nL69lGlqpdl9ymbRJ9tCBG6SnyU46URwI
cI0kbx59Ss3ugzfmPvVd+kXn2a6vKeVrDuVAjBRCOcKbHbUx02S6U394Aq3jmDxF
OjRQx/NvsYlje9Sl186pYCrPpM5QiZuHUMarblq+7/gLtT4FlbUl0VUqhd6gBCHm
hphRfYWARqZwjMYa9gU7QDCY96UhhBH4hvwYYdMZPJ3V85tVXzfvBreOBmnibtEw
YZx6FSQ+P058HwhLMLyOm5+N4qut/eWh51F/NVfbR6VOaghzk3IgWp9dWOzFD5rC
n/L5pIBrf4CtbqLyG/WviKYd0JckEQINh0uYOSonaTVThu2axwVqqdY4hIGAhzNR
rMO1Q3lrddwwF8WlRzboul92DvbpcwuZh+6JtwvJE+yWVz1TddsoepPdhWYRohY3
dDT1wwGBfm3Z/Mix89QZWH0nD6rTsfQlm8OkTzwgXXR2PYtbYWB326KLG6XuRfG3
VpBfTKTLWCa+aYe3wTW7s0+JhTd46xak2upMbKVhkg/NS67xvHxnPbJTtDzHrxPw
ZWoRDJNWipsMR7cssteBN9kxGuRks7fSgeJzy+Pyndzuvj856yJfnhgm41+puB5Q
KZeH1HkOeL6+xoKqxJtfo3INlcJXjAdIEs9PC+sKWNefiKVCU5bGHBsAyqfDLBCk
qBUU6mXuc3lce+bD8nSorv3i1Mppcla5M8RoLfGiW7oTKCercKZuiaaY+9HRQiKp
xNl0LfaWiEQ4QdQI+NrAaRDXYZL7lyH88bGCJjcQI4Awu/C3HDZ71hV6OQfo59yY
chp7BdrGOCH18sH6TIJh70zLNW/yQCDxcXHVZQIJD1Tj17OeUMIyEgN6u0Sgeuuu
k5THJZEUEyyUzbFZ/P2Cypa2pf2fP4PIaWSTcilnPXwA0iE+1EmXBlVYYhZZI6/z
Wj589RPWpiSHJsteGsLWcs5cTvacrTH7MPz+1ys6Dgu8tOlTZNkimW9RwwlxRSrA
+jPUU6szCD+gVoybnJod5I9OG9HXP3ZkZ14Gsg47zYHyIWKSLTH85eiP4zEPBtS8
UAKV8jB0+JYZc0oYhI4LXuQdtG+Z/eynBsffaMG/c/sDwlCLPbjmofCuEd5pDgsx
xC9nuToBwpncuBfINeclsPcTZdmVB4Uuzy2d9RKMFEGZn7LdcUoXNkQGVYOaqhh7
UTF8zJaHneskRkRQSC+IxWgnVLsuEE7inH+lQkHN6FGwUJfReebAeNnQy7lUp/7v
jzvWOvtBKzwkOvSbyxPCmPuN3KyKMA+0zdzeRhCSbnOST2WdVW+/n/r3Sc5a8EC9
uKWAEYZfOfCb1M7mmxTUTtr3giTuBjpG8Hbqd6U/H78Bxn0s8tgpTMUk8WlUxFDh
8b7+Adr3FnhEXqYkQipqbcR49hkh3lXKbI1nPyFzQ3IY4NjacCxznBEAZ1EjXlCw
OMZ7INAPlL1jw6zpyAUBRRcRoaR6kea42tKcmi+pkNaqWr4791e+Xg6jdPNqPw9i
9SZrgNqjnhm5+DXiYWC3LKYMDKQA7ZmjEzaCsW6iG7EMaCDMe49NzJp1xwApAMBr
ozrzu43uNK+NyIZr2AmH0+O4z5t1QGyhJs+YNvUrrLymzk93hYSNKiz8K/JTv2If
JBqBMF2S55+e7XO8/bShdtE5AVEKEt8ZIsF8qDZjPRwZ4Jdg+EEZu9hYoOtLiC1N
1w7iCoPPGZv/adRaYpUVPzv1c4uclsVUTX5dDPz4BllBPYpaXDELWHqGu6LZOe3D
y/NLx8nTaXCVZ8cfkqJK9SIbWhHwCYk1qzCvwFjTBmeplUpI1VcSS+Ip/Ga6jJNq
mS+0CPNxsz+TH5NHCCNawPGNEsk0Z41qkIXGgsmzNegyoWlTJez8g06dH6AoUDfk
lXpYgVAwtFW89jcsOhRT4nLH5OIJ+zbrbbIh5REtpHUVDLXaOtXWItbrkt2HHnp5
FlPkcusEJBS8QRxAeyjxP06e6xw4HibMthecX/CM7K2Qw0iSzEyIpKjIlCmuihfl
bevAJgFKRd9W5fS3JcO2ZqEZhLpU5F8OqZsZorrfu353JGJYyDD/c8wkutbfuISX
GB59HFxHcdqy6dszInu388O5Tnw08uWJD3i+9QItEYWqHOXbK1yXOGVxu9jb/x/4
s7FGzwbMqbDafsI/uK2tSaPaSGYv56e6eFYn3ZDh1+cRODJD9A0e1AnbaAm6y8G2
xqj3xjM3EarjOy3L8MMXyvYxjYVD9ddbKS0iA+HHtHuNmHHSJ9zqUIa+eKhHSNiV
7via2yIuWJmclrHkt0ZG7Uzj4Bvh+jXZ9UQT9FdIVaxPXvMw84oRc1I1fBgOYlDA
JzQwT94AoTtTPze3pG6YAsd0hlFiRZ1BZaUJmSHRdD8MWJmqDUbQThjZoFsly1Gj
UQwkDrkqUlzRjNhTOhyloOiJf5nYXjcrKV5+yw/iWZvH9MrGBf5jnaIs4EOftBkJ
OEul6V0AlhZ3KeOiHXmgmUaLasFZ6+yeIWN0cs0tAlSxlAucp6qwqx6NDmR2WjZM
hUDnfLU25LlctpluHPulZlaWHI1SD3ZQ0r5SHSCg0rA51o51d4Oh0SFEC7px9QWL
y9d3OGrs5I4itHe3AWJmfQdZuOaktBgyJNfBK73xWyl/6ckVnVG10uBRD9y1UOVM
U5dEE2DNMbm/Z+166BkPsdAgR73HoU34fiL3WH1YwC/NZzOiq5jCb7VnKmqHtwbw
OTktjUYugO36/AJluIVdlYDy1SSdwZE1WubeCVf9PLcsQNvOs6F6KNJp6efVRfcK
XNYtyxEAMQ5kc6eDum+6lFp/QlzIJumonnmC0FLymA2jYFwapnHzU04tlx6xURur
oXMIiwAmPG/bFZ28alfAo90RQyXZJ2sEfOFDBgLeiLNtK5FioAb3F8aRqGUbLvwK
9n3+sg2hJsK0Aom5e0wE9jaVp0GVQ3zDkaYTRayx6JKbTu9Y1M1VzFdFLIFIslDI
L+BRrA64XIHLIEE/hsy88vUDH469PNfRxjy+yGgCe8BwnnEmI6fYS4MfjD1Tb5fn
nXTAAhP2NUMYlquevxSSINpwmXKPLxsJHivlYS+WWVr1084hd/IqRlz4VU1P9HBc
1CItxOEua92YqX7rhCbs8XfYFImKrSqAkmSmLaP38G/kD87sMvL7GZfzh2BC5eUW
JpWot5y/OSs8S59tM4Fwm5kZ++h/01AMI2h+LuXSsQNdF3knuONWEaOzkhFAzwNx
F/LfhYhSWYF6U7ZvCcSI+ENqS5G7eqPpkF2CUv9RLsp+Uy6X5az70SZAyY15L8or
TM+egdWRDjUNpuF2GxeY3olhRLxP8ySrb+m+7hoYazPM88tD8SBnQHHF4AyIGqzC
w8AnlYKYygx81/FuSFjzoe6267d7ZFrMJc1K+N5bs/GwdfjF9pAMDOVzZzaGIsrr
6/fV6Y4HhhYOnNJbxzc5D5Q3vGEEeWAibf5apgb9Df8xZQVuJtHH1ilQqCGZGmbi
N6bks0ByJUJa+k177ecSg0hoOJ09Y1TfMlxkyGcit6aqLFDUINmb82LMvTUmxeop
Q/6xY0gj4wBvilcU9jQ5qBdHDPvwXRnxTap4pUtNQUm/RP+5S6gWrYEchEl77K0R
wg3AWoIE76+25zfJ5zVMJloBE/sIt11bjTook1zQr454c8LLvCVpFv4qFvF3crYy
ixtya5NuN5XeSbmxkslurZCSiukXzZ/4Ep6rVXI+POS9lre/yE8jFzi7DYZo22MP
hbY9i/VSN7sz71JxVP9G1OSHeymw8Q35GQ+LfLwD4iKbwZigKybTFAufwNiQ902c
zUE0apMJ/SGMldCPY9RPL3vxtcCpUgavgXLgZI7qUAQnSb/4zc65Syrp/L8LDNSf
i9vCawguTRsrl8qmFVrJ/NKeUQq9M8CQliL1gMX5UNZjDqj1+2Eg3W5ANczKPy2K
FXb/w96rrMudZA3lm5ilRtrqWGHwm3wUGYUlTermHpgaFoj7pDWcIIc7LCRS+VQT
zl9bCFmRGW6CIK2bqXxIujnJ+9RADzKRIKeGV5uyPZow6XFl70pLpw0bChErVdwB
uP2bza/+/lio+Hc09cyAIGcGDeFCMjzK4CDsRuRrVXZKhdilaNoFKV0G33tlUWJG
LqS6xprKlA3t21ilQq/yRYPsAaFkQrDBar4lQJMYkiyxvlgQ6FuH5R+mLrt3yxHA
OTxosBABQcHkGhbYv9z29o9I3KZcxMQ0gqxNp0HT/xszoamitJBxOM3FybX8QWzV
nl0L+zbFGmFR6w26Kc9fa+lYpIxc7Y9qZc7Riz/1tsqa87wIfU8+4FluoXcUi9wP
Q7TQbeYbnGmBU+xQlJmP3MPZ4GaxblPEvrwitfEjDF/IiNWAmAz4/xD/vqwwO8OG
phckegp8eussICjsD2+EpGeyhI2qI/BS/Oi3UStCC+I7kQVfxOc6zKUqKQ1Ou803
v2UAB7E2wUfrYWNqaE4o0BbQGRMiwFqHqAmtAOh9VEMmZe6ngZD3QZLoN3DVz2rY
510SlIq8MI2DGFjuZQlB5voPpa3xjU/zwJA4XCmIjDu3NCEjWzIDlkRUHtHbKs6D
JpHsjaWRTgV5IRpaU1SuWqhcIbqoFMhvPDF/kp1C90fAAb6nLIzfVKPl49ye/hJp
bPGAN5FzSDYF05f7sAJnILdQAOtU0rj1FCU3x1LbFjqw6VfJENv8cjkmdW68rrnB
R80qBOYAaaeDjbXPamgls56ssDTxRFI2JrBGdtllPkrEdYyfnENyW5Kl+n/G4gHQ
RqP/xop7hF0aYkzNmW/6HOlLr+Jn6/Gt9oF5A97uulXXNRojiaf3M+Q62vUXkuAa
+3uTe3W//9RxC9s6fzT2nRfkM1V1sB/wzT0CbAbyRLP5ZfU8pwulAeaCV4cjwKPv
AjvygUb0YXaP1Zl5zrqGhACTMFPqc6Pnzib8GFxnbEIljNBx3rdtQXGX5L4IoBUX
wZsFuJEWJG3b+x+Nq2sFOqz/sZhbt0qAx2tqLnGPjMitAu5AySiSzlWqB+b5jOMa
YRLNtzev/cokmsuoopFlpwvU1LNsBLz8tx9uBtWSOIDWJ+naZBWuYD4RPyhBq5i0
dBv/g84c9lT34Y3cRXsXbnngbjnXjed0DyxrgTK4Hc21FyN4XjZlWk+1kU5HR2u8
mvryin6JQ/OqFhrZ0658z/nIoOAUKNvqfHMeVlwTx6pc6iLZaMvSWDvw5u9tJfpK
0px5gCmsE7OasLQRcPM4iFDjCNGPXc/65uvQMZKnW4URnBKNu5ZszFtroIyB7LdL
MwcLJ2YMk2HtgSlBmJliaXRXEdY4+A4+jmy3jWju0XQIgcbyanzxS7IhOD1d694n
x0sihPj4qWBttKTq16G3O+eWcQZpVZGQEHyYoAladYG9dxq+Yjvq1pdxyGvHSNHu
0Q886zxLyCLn7Fdr2/+TvbPcDaTI+TwoAPZAUVsXQ4IYkuCnPxlrTlmcwQeRRrLh
gKeac4oFJCmAe5sZC19x83dpNokuBxn5Oz1sLuKe2GbMLK9MVD1i9/2AT01zCg1N
qjQph9+rETLBx8CHpsil1EHU+RVTe6ON9xs7xXPUs3EIayBQkjH1ay0VULHo8fki
v5bf8POHRD9+LwzwUVMXQI7mJEsRHp3aTtT9axG/6eCuNCsO0Nfi6rH1dqy7oTjt
TdidDv1O7tNRgwWNsqtifrGiyEwt3AnK90R3KJZAyFGg2jMZ0ePr8m47j4zfC0UL
GbPxP9dtxSwyyEu1QKzS6pFxZc49YrqwDiwp/HXRueU+K54QwRzdo+th1GwbzFMr
N1cZO1Afhn0Yga6DrKhF9KQ0+E+lz1lDAbcQRd94nU85sh/qNqD6E2Twefyg79VZ
rYlIaJEmHxabgxkQ1T7i1CmteT8DvjIlqBxTHWhNRJ0yDFiUjlYte+x1mjbbZUfN
oKuMsY8UsVGF09T1AO24f72O9rGOvKCEbFULA0+Kx4eaog3rnG0t1C6MYRcOWcM4
0FlgbPCBBYq4zNVSP51yMfa/vhSbXA4MU2p7+/bIG6eO9XTZimf3D647y9Qly8AR
0YVHPYfHuDvE4Y/7s/v4Q6IT6YsxBTdkH3BWSHfp6171MMTJkXn4w9eRD0lXW0sZ
Th22xJmK2z9IwSfDQEz+Ds5ydAeLKrx66YWgUyQA9T9oEka89JuiL3i1fEjODIro
VZz/GxBLPMCz2s911wBLJtM/ah+KxkUa3kznjYYxs2IQMnvLabGY+6z8SR/q4wGj
bzPvUzajWUVlVPtEi5M2UdNrlfnOxoiSk/6XyBhmaYq9Idj/FRY+X4QPqikYsar/
B4/NRU4LRuDW0qvd2fHBLIEz0MyvqiQZ+6DlrG1kmBA2Ahr8gCZUJ/iorIwlVUP8
XHvZe8+16PfbarHFiwBu/FMoRE9WFPlxh1GQv6GvlhAxHb9ZnfYqqNVi42fI6hSo
DU3FcLT+NrEHm3m8UJegxNnwCUFILdKBN+SnGBvP8sSaL4Gw2HGICSeVIGq9hdI5
luqxn95ZKiN03Hd7kdy+55rLWtDSAPzqgvkRp/0AlHYRFCpvqgd3VnPDZABVCvP8
YM34NuoRufW+8P1b4YnJXFm/W/bBumPS0QSAXxquoDiUe139dZYWysalzEu7yTdZ
OiKoQAfsoYYKsKp9P3Q/qalcBkHhV4a0O12T0eoNJyIdw3N4vF7W14uG5fwJ9XIA
lEZzA/PvMreQZ9td3d8u4FeLFm/1FO+WohiT3+n18Mggj5AHdPk9pAPz1/rrnyC0
b1s2wK8+3Nfe0/YpqMC8JGruyc2mlnd7GGJnO1S7ZhLiPb51BnPX8Wn3sB/1jNoa
A8TLB5qs7ARlTeTRLto3wNX6QKqmLzOS+ovKqM0MtTUViL+vuEjozqaCaW7gp5hb
/FQS/7kfMvv7dbm+Vh+ruYG+YN5UXVpbPiQ49IFv4R8QLmzpORDHQUdv0Poq6OYQ
7YUS/C1wIdK7FlD5a4o4hN49a0TV7R6PcuOngux0w9kdx69CnKBdHNqKr38jv4GS
fcMthDeXhReZg2/heUSIdxYRH+4Wc0f5pgyZwrN1lBtP4TVKO99nheeQledarWlZ
7JWyHTFOmvxBcT0EAInUkVPkb3SoQBKm5/4b6ELLsOS9OQF+47tUFQt9QP5tYZnT
JfdIaUqDw6D5G2PksQy8zo1F+oMkgfSVRsA6WPWoKOENhHt92FiryLti+ema85Jr
THjBuzj1rqKUMFuK7h113PEjb3PbbDaFvZUP5iCOJYarNS5gctk8rfUOA9soWhJC
ccVwAljI9CbFcqvEYSf+MXKBrtb6JODV+lBB9jRsXt+64OKnuIxY5SlS0wTXiucj
8FuKoxhPv3J2dTGI7seg7XHMGaK4UKSjsWBkElxthWTFh4cECLsWN7uK16IbZ9k9
4h3aI+CM8sZ2l2A1Y4vhxubm2N2s6FI7kKFrsGUhYrtNGsoAKv+6nLuMnvR1GSli
hs4iw5QzI1TMKa5IcTSGkLuOqmaF7KVuF08wmE3cySMS1lho7OQOplFoN2OSl2Hc
RxxIBzU/UH2wPXqQEIJ9fKqXW3LQ3K1jstxTy4d90ZG1o8kgb4KzkQ6ZASgsPSw8
d0y4H8VeDCIhICs+Luq4jUhFT6OkBUxlFm7P4PM3NjkaipWBUt5peTAsZIiacU8C
iCFlE024VK0L3MgJhkASVUpDfBzz19ICoZzsP2s2uNUXfF7lZwQBUJ3yk3L+tIc8
PJbtCzty49VRcJKvoiluqgqxFtBeYWtVJCnXVbi7jbZ/trbSdrvwbWG4XpIKV0VQ
MvEMw/aojgWjGJdofNQuEt2gD4oBXoaqG8lY3zEhqW9FkmOq4L8PNwlQ5iSNhdL5
9K3/iTBDPL+x73oc+t/idiQiLL/eM0xq5fugRLMce5XaFeIda5bUL5WpkiZp1PPH
oGbcAHdt4Uaty96D8cRWlkw5VWuU00FkvRTl252t1gE5ouI4Yz7K/zYR8Xkl/0dY
naaRyq6d+tFYKeCx7LmZjnZ/oPJDMLIfIeixGGomMZmGXm+iuilr6eRiZqzHCK7t
U/XSmNdA0+kH+WU9BkDxLDkWaNlJYyX/UQlOt0+VKqAFKvxgXPm5HUED0U5Fjizh
au01ZaTuestdzKFe0sO6cERQB2IEPAieNolqdzTLehcWQcjhII4xzTw+I/rF/PGV
kbibKx8P+xDgFNxVVqoR7fgbrvRgGuD0oLlnnZl0s7dUnZHTIhSWcVjJbEeS3gSW
noGKGIF6jPZawZPAidjufs7X/jnfcIKnzWC/KYVND9cbeOADPabMFsKcEQnYdXhV
eCMuq751P79DLfBFsmqkJj/MIx5+L9gi7ahcRlXiXaxG1hLoEohFadw68HMlpf3j
3Bfw4omhQ9CxqrCZTVOV6OyynILtMS5gDWBpNmUSu4bzpBJGV4y6i03G+JcXtrfl
6nH5IGnaD/UGElcxYAa74hoX/hH2k6k6wNslNiuee8411PlyBeLgGetvLhvI/Env
uO2oSxZj94OkqETfAVzNSZhOEUJ0kSPVysB4nx1yEGSwNaSd+NdH2WsuvV0DfE41
n23a8P0hrTZZ2Q5qEsMsiPGx/tJCIhhsrOWwoRj2SnW8YqKppOqJnrhhFmISBzu2
7ZItjJYu0NFR2/czdDFbFbZhoQZnw/VvidFqTpX7HRbJku5D1IrJl/pnxJAU8RjQ
fjRD7Y9NzFl/nl4T9szQpg+Y3Eaz9s6IGz5AzGi0U0q7a0sqGFZZV+dSC2KDZK1j
sw6EaQluk4rIWClJkCEBzC9D21uo4jtbb/Fba8okaTs4ama1RI2ElO81qpzZF2Tb
pVTjXNWrR4+iThA8PNQJKYO2ra35kcSbRNfTt410ai6HMdRn6RYI8FTj2m3Mk20+
dgag7KN8VAOw0j66CrRHOE3IJi/gw8uu9pqqEf8nrSsSg7I7Fr4+qxQCSf0sXTts
PmevWi2LhCbEc8Y4Gz8UGL8kW/wgp9iraFT6u6Gn6EuNNd8w6euWK424DOtR86ES
Wlf8UI2vNNuoK3hkmxnbGllV6i6IItW366+jQaYgjzuk/zQDQ/EjW+dnblJ3gHdZ
V4RIJT2SUcJ9FiG9F28+84U151Gzk7EE+6+5/1G4h31EUzcpQNiLXYMv/dnbtWUU
L3Pl880bTfN9tFW0SzziLOOS64q8tjRqwqOZBcgJks8RxmfGQNr2pNXBAVoelMRW
FnspFICOpGTaO5XCkKzcAiQeFPo4Hj4VMjyRWmWoi9UtmOW+luDGzC02aE+a7HPf
M2Aygt5A3PtaawIbHlTy6iWK7wT2P2gFfh2zlTNoXG9d3UjqKFNeTchfHrvTUCQC
1/Am41RedDyX+lion5thA+3cO/eUGP2sP+B6LwvLSAvCym5Ob04cerewQBXxNCdQ
hZOQ1WPNIwf/Ey49KO05Sc9eFKBJ9Ow05bVe2HNitpK73TMbtIILyM3pROXRCBpO
oZA9k1/5WNE7gSqoUnaruj+D73dviejcTvODGr0B/E4OZwFdhukCyBErtidG1WJy
DoYacaG4UZyatuYEXg2jTV1yJSzVJvQq46qSUHwAjAEUdREOJa0XGwWu0k/z5J4m
c6UvnEAxsO46HrkTWnSWoihIQm7AF/uLnnLVL/wAhXsCDk6q3RycYXgUoSh1YAWO
U0MuQ3FfoAK9pn3P3rQlPPu+GjBQaaA7pIVKcrwV5bU/JNBDTffwjm3KcxUyPI+l
OcEsMcAVoxIYj8bUROQ6cbaUStWVGtBGLW68V63X2hp5JyCzsKuI5l57bCEmobSz
OkdJZ5nC09RQTfD7vKXapQPslmawkYGpAzYpNevj01pgg0GdFnF64KJUljN18K02
wRzoZPf9pGKLlFKBDczB0w7irDCjGwzp1YHhSq3yiX9CSdHqDNkSXkiH+4pAtBnC
5bEqE4etT9ZUrWU+o7yvdyRIM+o2qOW7uOMx/LBMaxKKmuOQFXOxcYWWTTjjLuPj
aAyOYRbjc9uSYu+mFSzk+WwSZwfX0JBI0rOaf8K0QcO/LvQnDIS7DVlDoFmJEstN
5wgJGP04Kq37Iiavxo7hbO+SXZf4Nigi4BaDVMvn2w+i1u1g9158UQmw7/Mkf3ev
KYylWrSjOYV0vpBjk0lMeNf5k8WAVRqoHkhuyetJWym0A1mP3oqx9o2svWEiIynw
ECRaSb8T5jb4ybTZesQwm+icprr7ZzGZoSYxsryYisoTywK4mhb2rIhk3kePDfSz
LBTEQHFNm/4yqtvHIE39yQ7SrKtwnfB14M2l1C1EWkYXNOuvEhXGdz4W7qZdoOCQ
ghxJFQ978xMktS9B+cXJtvgjIvpO6RhvZcrfIwg7uT4gaCcWRxN/vzxKsyQw7HZ7
edr7K4CQYrZzT4dRvWh6/hIfVoiThwLEgASy717aObGXjlxGPqZz8oXhwHOqkC0B
+Qw6cZ+XyW4iKsYw0al+D4dsFRGl/3bNkzStK8zraXvzdeXCx/62CooU9zZxOqrD
ArdY2M9kbGSv7Fu+GnXMaoU8Wsv5xduMlZDAAEz3BecH0/Kr3EdjaxznnE1c1/14
FLvKDSFOddNhmIJHIViT4XFbjT+Nd3ATdj3akf41vxqkxxPvo5p+S0pcJpKSBFXd
EdR0cCU87Ik84OlLPUd80f/H9b+gK1N4SVPDGzFOq37zZYSSrImoFZcn4XPAx2e0
cGyS9BvlMvadZGpzSjDmXO9uhI4jenyPiQGCIuI4h8E+vv2ia3uRX0TWYpnMkTy7
x5ByUjsjy/DDDEWP6gZuFdXUbLJjMNePQTb0M2SZnSvfX4BrtmBrTMXY7Z2dK3zU
PPRBRyvbYIWBgiXsMe1sX9Xwt4V6WO8BquhmfYBPUTk60xSvyQmBlXgc4LAxRyt7
wt4Se+7jhENF7h7wa+B+t4Wc1xnkq4AoCXUbBuV/jF6q+0wNt5rli/KZncqexFOa
kA4R5jBDRi8XjYbY1+n4lWk1RfGtVqgry3YRwbcGdbZkp70CAt8rKTM0tU67sGIo
5p2vEIwQMiokvLZH8TUJll3xDFJyT45Diz/k7M0EdzRJxdjqKBebjNlw19UAR5gU
GgvnBPv0/IWR86d1WV6S9WDjEsIiaWj20iaM+1eydnzm8Urd6wiziqpSov5zdCdn
dC0KIQ3L6+AC/b12NWnRS8sJhtjUgK5BRi8DaiKIc4kUnLXgUG9vWwtKBE5Lk/Lm
etpPZQd+TzATFVqQnaiQPw4HkTTXR0SRJa4czim+MICJLDhNEQddIsyWx6A8pRK+
Vi19bFQd4BNSxovr3Ell0sz7zP5W+DsQIGz+UUyHK4MnxT/S/B+d2Ti7i2/MDkYJ
1WrukdtEhcTg43jeDe2zt90n9Atl0MI3D0u/vNuDJ7VQImvyGXuPeUO+MiCn/gAb
ot3FVIwI8CavQYdnrxrdzST915e4P40HxgPedvQ/xI/DEAa9uJ9HhZAI8OQyGpE9
Mah7nDhV1wDRsXz8yksO2TlBn8E1jOcIkPZzDOvprxKgjcuAYPYynuNjQIico/F2
wFnvOS2N8PFNfgEiQuGAH1+Oc9xDa3G38/lL7HVsAX1eWyAujXs3/kyLzHkgS0Jx
x9TDxNaB0/BTRXMEJKzV8K/wjwbHsaKEWT7Teg8Wo/oLiHm6mHT6mKdqN5xgWh5b
LxQDKonxzYLDUT6nB4eQluskOyttGCjWqCzpldHb4U9WAwODt48rgkxm4FRvv20C
rM80N2PTvST6ebA972GCa4iT95LOwnpYC7EpRc3DUk/h8vzjNCerkrvSaV08axQC
Pq+wYygcXbJP/Gk9fEa6w7Rht1pPR8B/R0r6t76qYdUmEZedEU3pw7FNOu7fpKTW
PntH7/cHvA89AEvPL3exJ95uDN3dXKQb+m/9Aj5USjVIS0aoi4IH7703fwmLXpLq
P29smk22hEpya4sE4o4SdvbKynaUMF6wlU8NX31UYGpWFcsjcSAozgVS8Un8Z7yf
9KWnNfse0CCsjBPSWFUT3bhNerE20WmfsLvTXY7u+4ekbD2EvdEW60sd1luP016Z
Ryf+m7K8uAlTwLiqQiQsWh6mUFKihwd09KHLKY+mj9B+k0Fxuq5F63iQW9ItWloy
pTW0pUWlU+ttkWoBtlglNWRDdG+RZ0YCKeolE9hg3uFM458+n1P4L2WhMuSMmWW8
rq/O4lyUEfttyCnHmLhkJbMLgghmT6VLcdb8ICCEM6tyiEEek7oZxSiVkvx6g7tV
wkJlPqcOLrYCdhlRlTSvyVpY3PhxXu0x+mhKig7bPf8186PgXa9x9eBS0z1j4HkK
mDxMXk4qt2xZkcxWq0ElgDdOWufTBIvnaEWNRSq22zb+iSIDdAnkhtxDoyleGHl2
hCFNIsUIeGzlwwaI1UHGSg9VDOg270GuQrO/F67TLRP8Rz6qpnLuYVNroUhoqVi6
FqUlwIzFDWmRBagSMZR4wYkvuD6E4YVLNSccSgqfnUtxUcQsNACSxUxNvR0DjwMW
qAAAifdPHVL/xf3hV4pVa0Um1q9aRbUYd9mxft7CSKv6Xdzzc8xLYHG2RDLZZtyU
KS1G5bu3IBtFTrsuFiafOaUWSrC45k9anitot0MHLgRUb0U72nY0qeEOVluSek9O
Ieypcq59U51BtUrOoGIJd6KCV/N5z9kikiQbNd/B06A=
`pragma protect end_protected
