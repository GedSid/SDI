// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:38 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sHJWhbZiKjSZxz+LS6HaxJicuH+rEVnzPLlqhIOokDCZtAKr7REucqDREBJX2woX
ByBwWhz7Mx6P/88bFh6TcXKFsNo54GnZ5N4SuIryZMrDwODJ0q5N4Znf5mlGWUaA
dagOUKkIh/ZZIPErODQa1ybTZ8J4IWTucRtOEayM/bg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10272)
AcyRgLM3GA3/m79ue4lYwiaRyGA2ZMNIrXx7lue3p5bwmA9+mBk0nwhTNRoBx5gi
c01zV6i40fJkcv8nSAuStCBmCFsfl261YLRHjzv21+n9+VPN6YLnIxBgqHrKZNVT
FjqKjfgjUUPYt01nKtHSD27MAe6nL97ZsHBA3JVq4GiZG5lOm+OgJRltZIyLfJEN
oPW2wGzU40YUtfDL6IL9vWvv01lywOS8yovrHiqbYwZuPSLMLsJXbyS3rhGTBGov
rc5DMXhOPUH59mEm1E/sgKTQm23a0qmYZYWRoEnPak9jXcwZOaHpoLJS2Xxdym4j
V1dzlZC3B6n/QMhA8NC81mJ3GP7/TW1XNv5nnPtExlLSPA93CsPf+vKAHzXLdSIq
/+JDCHBACE7/nlKo5SjpF5pjVAKhGYaXblR/25+OyayZ26r+UhOlRmapDR8fXVdL
QnK+BBWIhKnb86q7a/E4G0u+Jsio43pVibN3+bl6dzUcHTOKcV+4iiwxG3dzR+LC
5MwKzX+d/vFzLSwJot/X4ZKzdESqPwMIZYkpMuPdLm/LeWDEYEd9IjbyzLMnfsaB
z2SItzcNuB5F/NCj6sCBzBQiRM3eI4e1R9DDaPL7WB9GIgaZYYpaUPlvBrQSXQ+u
B+cu0XV5ml2afQyVgs5uIUKG9Hjk7clIhf+ESyLxIRB+7wEDu1Rcn6PYHl3SggTc
BmRKknPtArktpABTQp4sztr7qZhhkHO0ctCmscs7xmyIeYYMd7oSVk7XPcwjSAKW
sUw/fsvCGugupKhv5UUMO/z1M3eD7Odn6k1noXq39mhcG1ls5J5gOUHK/uxTQdB4
JNvF+ilTCBQl+QXCRz/TSI6y4HEVZTF7IlCO5bPn9PxBlA+jivTK2R6igKuCDFsV
L01Sg1T2LpDZdXHSro+iHV+T02Q+6//4oCS7E9ES0okX1J847ySGCU//IXF+ovKV
PBQt7jv7Ln07zqdTbdkh0sVXopLxPvti0JxcB5uF/3G9qU+C3wtCrYjBe82967tt
7paotUnZuCVXyglT/YVQGL/qdMTWNrDJdArhOsyPg+SP98nEzJL/eovCZHLcAAy3
8+xzkO8I9k+DvHsdk2QyEe1VyDAoZRWroteAtyEFA5lDiQK7rBwl5Kw9wVK1UFKR
j+rAFDeyxoaL4e4GwS+TwFxt63XTw/cpw5DhTdF1+72kzYHDJe5qTzoG1AYnWwWI
q5ZYJSmJx+4VR+cb9YEYuQSE8/+/GBbG0jbacZiDPzgEUHwb/XcO78AxecTXzvKr
bxbit6XaveC8f8wW/zpHL3fIHdp/LEjnlZsU4l8cVtphPczYoym26crCBHVETAgc
UKiNTi+nZVvYCw87ANlRWnUliJkM4ZxczzEXqqttNAK2QmeDeu/VqVZzPjbaCsjs
mLgbmv0WNPDEBvqekb6fnMLhiCpmCJiMSNems40IEfbZg3KUercgm2Padu0ncmaM
hEwOkgV5Ckua8lMRf5DseA1ck+wmpB7lwThYejWNrrsGn5rLmBk5idZy5p3T4DQa
aOCI1+9YWPxz1a/x6LLk/bqmiqKkHKdn//fSh76dZb7gTrsEKooVDrL7c0pZaXu2
8eD/qqwQz5W0JXmP8v01TIbKUYOlNAgZJ1kNNrbKB9wxu/a/A9NZLbJDdLy/q1o/
OUdpgJzPVsDwWZPjVTgcjvHB2k0t8w4wKgeKWQiLXOBHdQQlRb9+7oAaewjUSOgh
E9Q+ka/Gyd3/HC+XJouAO2ktjgcWHNUyVvEbvtLjNI0vG9wGv3+IeyUatvRPKzoq
1Nxju975qu9MmGL8PNja7Bmtjw55oSX0+C0YYjIecTeVKeXduBxqV/6Xf90f8CI4
G9nJSNDQ7A8xl7MAxcSpSBO0M4Soa90TNJm+JxRJLjV8QsdAMBpsgHtizG4rUT0I
wv5M9OGz29NjSR8KzXm9DP0inlQ4m3pwdsCkixGqvn8IxIyEWDKeK0PNZB5DrIlH
VJ1VTjh9EpVS9QMbSIy7l/tYmOxUCEZhd2MLW5ShOds4yGje/RP1Y3h1kIFKNDHL
x2VlsIID31CqRpTXaoJYTbIg+W6kt6FIxwMRwvTOTj2/JqvGxOdFQ+skalReSic+
cJDtvy8U/CB/gbXIDYBjxgizoeZI6nbSBySCr2jSj3oHyhx2fo2xbeFZEaH01meC
UFKJ5hK3aBpCBxhz+Cs6R6u3asYMJr0nwt6jFf79SiUEKX+WLrajGCGFX6kUqtPr
iO/ELgUvgRyRtxAVu7NkUrp3d6NxSVjRkgwk2iHmfDu9iQvaxs0cdzgkdEhswR4A
4iYBHD2vFQUgxvczRGOe+DkGSlAiKHlnLakmGxtRjZjD1TNf9a/TxzJq0F9UyI6s
560f6Gbm0Ef6WVNBIFAaEck5EeaSQl+MNBUifobu8Ir3IMF2wU4U2u3t8r8I+mNR
Cf8V3OWKkLCZQrfjMC4Gnzfd6zDZjbV4wBAHOL0i3FvnL440d/hNjlCz11VmhEM9
Sy4GG16FoMNlssMgZ5VPKXM7TS+VDCTOTr+bWi/BFyKrCTem9GpdA5SBYMOVTZMa
8Ae6Cr7oOWCbc2hhzrV2fwE4yLuGCLkGH7P4hyzf2zmjS5tIhsGwAeCsaVxj55Zl
rN17WuyKzfaYSsk/eUbLoJ3AZmbEOU8V1Udrvv1EFHyc3a8/LIK+bEbXZ8fvGQ3J
cr3UkOhlYR13katiU/e7tH0xacW7xsZ3p0vwa1NhDzZTxfzkrZTQqKFaRPCQXBfJ
mNf7uPIC5HfIXU7lZwWSUhEoPiwnpgnuR3dpDugJA+pDDTOgbH0Zm0JPUMdvCQE/
uPmlaQp1ArPtlgWMWWj5H9KV3CbUAzMCYYvNFjZD8SftNLesysFIFkxXJF0g4zuw
6vBNIrgHNwuCcVX5Om/OyOomyIaxIheu5B6j4jPJtvOn2OWmIwP8/1gC4qiG99y1
k0bYlUGvSMZp6uWRP6UN3Lc3QuOHMpm0PBcGXPxj4pacUgXF7uB/HCRqAGr6pvPv
oA64UrYpz44sydDbZvuLMADXYU4beicbPKGOz5cdpFGDBkBT9n/mtNOoNRJpXN3K
FJoS6QOp7vhNcvHU2K5TOZCfTRj9+23aQrK0v+U5YyyjEJJz9Z4YX0MD3SR6L7rr
aVM5kjUy2dHbBjBOpbk3c4gXai1n99Po1Ayhv2m+8qA4UV29fO5pZXdpDi01AczT
Bc/E7mieJJpp6USBkFeM6yRQxr4/FLkR77iLe18IwzE5JGQGp9k+36qu6dD/JmfN
09dXvEynPB8NUhxYNQhGuxXmW7Apu3yz+VqMiC+sUjUiQliZqGmVrbWdoW5+s9y+
/x3LDJnzHb5e1YhoZONklHcb4HHW5lek74wO0xj4SJgIixQtsgl5Sksn52rAKwFf
lYBGPFEqOENeA2uSzXiqtuWoKO3U8Abwrm+sTmJk7ZR6Em+Ig5pjZ3BAE60fOUQQ
2d9zIG6z3ZvfSYJMDcz7nK6MC6fFDP29ecmJsAM5ACV+Ceka8sVgydCGSbFJ8okR
mWX8DsSAAwBFb6cf7TLJwroCcqgQXko+FA6lUT1dC1z7P6iIdQsdssrHuI05HTFc
bkZoCJtyv2XnWE05gbrugGbpWud0zqn6h/cRrI1Np/IOZanOvYW/oeQ57HfPWTif
FwcJtNfMbSArfchaWjlf9AFBs7iBVCaNdwXnfab5MW1J2IcrK3/D1f6hJw+wHnJ1
O0951JPpnmC9JXAVSVCfHBWrxbbFHzJQ6fLB+ZGuckYLvq9c5Fw43Y+eAkPcXWiK
VjWq7ev8f0zNVx/HxJczLUozI6YfbTKj81rewHfq3ADPaWHm98QZfW2b1cX59NsK
kIZQHwbBPMrPOzrzqxYefht7tV7nPT9QhVPh8LG3eXJjHmzlW1wfTjU+2D1kgKks
VflkPcxnB0QRkmeyyYdez/XpkGuatDCKe4ZmAqWR8Hkh06h6jcWjAxEuciuJK+Pi
6KZw2Q2gOl6r7PfI1OghSZ28ek0mo24UNs2iIyfZhLeJ4bw0KEZTzcdM0kYpde8E
qeD35lL9Xi3AeXiHS1+wgyWjrlFHxFcNjQkmbA40HvnPu0wGoSyaMtosT3C8fPOB
5mt8ftAfPvNeYis8SSHeX9Uil+69w0Y08sAvtCUXPYrE3tuqBh9F41CLRmbt0qH9
LSQ0R0f9rHQFdtrB0fQEL0wHazAO/ncM1Gu2D3R94q5QrfQMMXWjQOXIpK8m2ULR
b0o/qAvrXETe16ToJXbYftmH+foATV/kZVrV1yHHbf6BSex6bh7TmPrgZlNUs3To
7HqdeD+vQBVLG6TrfRETVCL9KiYTcSlPCdvjj8QaCVuzUy0oS3/0zaIkfadRT4O0
23jsQEUnOzHlB0X916Gap24WYrCyi/y6CWAarJwIRMnvfdHt+V4eGAXQ3Dj/mIeo
8THQ9Wo/N+69IQLZr5pkcv3bVq9Nbr+J3uYymmzEb1lf3lB++fC/MQlUfwR2j4x8
S7d2PQz5c0oa3cqcirp+olQbeD5byIiJK1jr0XXPVfoT4z0FwlxpAzo/I+Hbm0q/
isYa3lWRO/GmZxd5AEOm0IfvRVwFoyTMIHSQOeaug9xKmyrett1NTHQR3D6nrN5d
o8ODWjVIIkhG2gtNZR2bLDzM9ww22WvI3fl2vab6s7s7p+9zYs+7AcPUQAHCVuee
8o9XAn+pu5QC6k9I4UmtN2HdUNLB1ttp3JgotWZphAADJlvLRvjEIgix5nqki4Et
1hpmIK4FjyOevxJnpW1dlTXL/XZAvw07smzJDKpC8w1W6KkI1Tf0nb0GYMakAmBy
PBJP60T6aYdlenlDCmNZf9Mhm4YhRvDsW59dgvaT73GjcDgiLiuhiNA5dDIgSSrb
uUs8MVRwY7bHYIX5hmf/Hh4vwXTOnMFvPkOg9yXvpIm5pQW8/NM8JLCi2RJfVXdU
+PNQ0dED7EvywthrdZb0nTdX5Qt8epPoEB6Ac/+zEPy6oVDrLDF6YyAKQ4mUvRy3
h3fsQFDbk3A8a7Jamwba3hZrugx/tKOn46thMqAHONyc2eilXKzNLrh2YsUBLAP/
LRbmjV+njuGkr4r2NsvXzO0PyPygwf/innm3wWGymtDRV0vsVyZ6O/Aod3lz/7mV
Asm60n0+FHPF0ZPjh+KH4svQS4J1XRYHl4Uw5mDM91qdtTY8A/N/AWgY++QhyFNH
3U65qzocTFICISESZtAH3pf1mUKUazkzqwQBIbrXHwBoNGlSyHbEiDlbQW5m9fNb
ibHxcytgkHLnvt4yk9fLoa3tLUNIiNV5ql6ygYsLFl9E5Kkog4B34ANDTP0Zb1sQ
v4oBXnrh0EaQE49nP02qOLxgqX7Q2yB3J9vBUuqhutwrZIZwmSLKjN3llPifd6eK
GNbFBIwfJ6lIKp+7avKNf9cGjcen65f7he7gCnU40VE/RNdcVBLFCl120b4ivVCz
YeX8FV4Y9hjQ4tl/qFyvHxA8bjTuRFnAvj39btpHHhvFJkS0HNNFrT94BRIrJ9Kk
nGmWQ2rijGgVcScmuu5w5ydEFZgmQJsU+6Mdh5a8akK+Ucz4sQD73DP0u5sf7Icy
mbkMfOffqe6zwYo7/o8tjqByNbaXAyyBAY9yMoOkZ4UG/cvR+5HgS1WYMitZQGEt
pn50aO05kjdCSEWjgu8fF26OWCbjHRm3NCvNSGBRPqyNFNXVS+I7ehdBYQlGCjmH
stKgZcEgAuBsenXUbzY0QedUdc331XgcluhncHD4KhCAPwu5UaLTPFd1QzUZr3Wv
vXrXOZZm7zEwv94uoDl9o9gVL4bZi27cB3DusTajdbjEoHHkNIIDiqtVpugg3tjP
sPL9YODOHUOhd6Kb9MhBmzXRJgoJOsGIQ/rJDN4TASZxRzBctet5r44VubnQQyTj
Q+Y3y1s9hNi4cJgM8rHfFef24mj1iAuWKL0RT0R3b40oeS8eI5MmhvsTAXlqnUCU
xD7QDZtp1bA2W8gXAXm9sDXBJxDWVitTKppcyqODfzFVN+1SnHXjDtryGmw+AcZe
3Qk524k9V+1smQ9xgBdVrAEyo23+mWxZjmHqjAm3ky8Zf/Wrpl7FDQqYen3dSeH9
tBsTpE+xGLkLY+s2lXVLhugf+QsO2Pz5UIHkM1N9wHGcdGRHF4+e1qT4GOagQI8+
5K/odHotvZpRDFaA32a693/n01uhdkUtMVp7xITH5t1eGWwdeeBZEM8HIqyVYkRc
IV8k+xse+K2i50Kf37utW4EB4pldSDZ026vDpJrHXwn/FaMBj0IMzXK4N8AQ6pRp
kOnnP9m9eEGGWAPbVBmm502ABuUkTRVuRyfGQ2hwXjEn+OCwM75L6UYa1isefCrQ
TOiit+1lJ7EBl5sGmIv+xrAyz8CEhNJMWELy/6moxtxnNx6UckEDErlmrNcgJyys
cnuqEXRw39B2K0ygf+nfRq6tltB6JPxEgv8mS9Q2Ly0jpnryPIbkItRNIKOgecfi
WMe4txs7NORnjngxk050qjBjZUetr2EdCrOqtXk7m/kxZrazgIYfKoPFMXeA6TRn
Lm55lzQSPGY7BTGF2sFMfpczwPR5+Ik+dNBiRmGOYM/OEhnszSX54iYmIqWDCa+v
xHKE+JJ+lK3LQ5SmFJnwwQq6gICSvO+GdSWGK379hRrgzGZX+2uEJTH9LFzM/zoi
XXn+Ujzjc2e7FEFu361VfovPNClCxc0YD2FQhhEBJlC3xa6nDgdVtTFw4UfjFXyi
j+mzmB6dtvzWKI+cIWFjm6OnKQp40Hv5iZVPP16kc8mY79Rgol97RdIG5ia8mXl2
v1uLv4p5b6F2QzXLXNMDKlway7PUxh1UaZExf0b5Lk1VkbBZvb61KaSwLuzteFNa
UhsH9lqC4RHHBWOa3II2sT3JOvdVuahWCV9IGdiG/uGQwfaQsxykYoh5zmw+aaA/
twbl+i3rg7JCXU5bwOcfWU4n/erBILfYwLuGjCEn8ijFPp7GC2OkL9gbj73tH+qs
fIVtCgUYJFDQ0jf2Nb9cfhxklscg7k3RbUwxyEIszccDjP0C4guoSoL+0f0g19Ka
+BDKQHKxqLyep8xL6E/Mk9To2CYZhq/rVRIJ1J1oQNRr2rzFvelyMd7rn7XoYK2l
N/czn0bpN7SR443tYisDzReR4YWcyRY546zwO2IipMRAaRdch9J02lnkMdqN+ZI8
038HqDg4vUEG+mGbCB/0uA5PjaKA70emeS1ddIjNsKkbCsLXudYVtGrtbIsCJogn
3Cejj36qrFA1T131W5OADgZZ6v7NwvgfN4me5gfEw9XM5EJHeRb2Kiz7KIH9uN3U
YpmOb3IZedvrtMjGJuyfgQhk0FAWlK4pH5HQt6uVGhkqQhFH7flL7JkUviqrhtMy
zT4G+P/h3GuokK07K6WVgHpa9nUaUCC9grquW+DADtZLczxr6Mv6kpZ2kqbfzGzR
w75hHUDiAtQK4RFBp3LHZNZPQeOoEsKR8sVTw27d/5KQaKd1ubkFdaz0C3v04xyf
wJcWrHubGqeQ5th1yOQ8fRvGfcVcqFr4oRvl4ynHLWPpXbrstostSGBS4Wrw8aij
fR4LE0OxGym7CdZvmg9VRszhuZQ8574ZT8OSr6Dwixr+p4/eqt5bWJd9aQEYxFue
cRzk11carjuTE8ZgcaZARVZnn9XC1kbJoxYc6cOXBag5WFWfBl/TvIFfuEK2sVFu
8bbJlez75NCq3gM+qi72YzUf/5T7jeT42RMyx+fG3d69cuD5ITOst8q3KmHQRb8Y
jTEvb5WNLgmnHDfh5ITNeGn3SC1vW1zMCym7tO99lz8bMzZ0VP/i4ArIDFr8d2pY
7ss7ry4vQ4tBF08/xFwZqGOiLUztHfGAK9CZI7f80+BtCKfQHw25QXrgX7H0doop
OU2RkilHzcTlqwRV7T2/XeKred1xFy4MrL9UREXpte9D+M7aCRO5cpZ7XEc0lYEj
R37c0nx4R+A10zrA7FtLWbIYMgOfpk3zf+ghC8jY7JDD1O4Jb44WJfWhyKKVRR/+
JBGF+1GyhGxsWGcmmLMAJQaRzd8I/L7Bwnm6NG72c0bmmtlnmdSYEhOCmm7wlNyZ
YMSdd/OCLrrGMirxrSyYpWH+sR0O+ZXMkAhIRAwxXniZrKQgDgBKK4gUZ4+Lme6f
kQotEl+A71bLKmB1quhw97PXJCOlHM9G1jKChyRJbCi8LpYuzQzpJ+VUGc/IkUsZ
+suPkuk+EyASo5WQPHC/zhG2hf0PeGNif/7H432fKIUYOj/AFIzyHxTyl39aHkvp
fMcY2P9QSCW+6/EeJoZZewozScHgoszCmfKKuhUpsT5xU99Hu5ZlRAKQSaq8v5Zl
Js2MdFbKazA8je0mw1yodXOH2ktgHayKDHSCnMh4AtnTAMRMoKy/DdAplQRnEmGV
N7MGE8EjsZpt7l2mOqvRytaGXpF8Je3Oa4aOkfJEADpVsgxcV1GtTsvG4ApnwYZt
b3FZ0KI09OFnl0+XzFa3AxgOn9CSn96ukS+uFdtx7wG+Bt1zfQg1mC9SuRMDqUgc
i11Ih55IoavLOqeaTZ7MMm2U5dH+lJghW0YHwPucctUTLOjg8E/meSGeckCrf88E
NWByZeECBJH/WlghCCnmcnRnvXH19+w0hOtz2uiJLP1XBLucVQQn3Rbx/kkb4FNt
0prvpjGzyJ/OzyLPJkLrw1PlCrDwqo8iacLbWLayz6ykmTyIUuaGdo4mY+SS5lFa
ImNcKGDUf+TIK6eOYoPWMooOTf89ebVyaZQ+FbrOUe1obLTgKcMlWSx7Te/V6GzU
vebM1N/p5ht92odUR4Un3+DVvtvZIpimv5bd3t1cioI96TjjX9TC+1Ty44kfe8gK
dYSPPnRwlTwJ5cfuKAhHod4PSRpMT0LUjAvgAgnOPSWqvCgSD26LF0QCK75UfY8/
x/WPogdUvcddzC/S3QvdSpa6HIROV9W7Qiu5PW7y8gjjyQTyC9V/qV0C4N1CdSt8
jOF/19jc6Xes6FiN3ma6Pv1lCRfiC2JXU41VFoOTn+qlVfy+vXAf3Wtn7zydMD7d
Bk8BiQAsSMaxWDMe29FA77lUi4yIe9I8nz0Sm6CYl855K1MyPOb2RCHnBsG87Sio
Ed+QulYTvkzWb94TZ+GpN0NliTHfk82Pwy51vD8k0i/vXq09A2mbje1MtSbTzAe/
fCSP3xL8YRMjW+EuXug4CrZr1dG1DsVxm9j+CtMA8O4gzlY9PoO0+RFekX0UvRnN
c+asrSnd2t3GRfc+2JVFA79HoX+flnsfniV6NjMNuOJqSiX5iW9jrjPD8fhFDGHM
5S6uChRjFsFg9XqwkIzadQosAkgifh55QTo6MMQR9SjIF6wO7DmEjPvVlQVURLVP
8G97NBDk2ZhYeTf2RFgbIiESMl+j7hOBd4xNJ2nQ8FpPLBtHHpHFcUECHNUyEMcj
m7ZmGdql7xHFmC1WwJ97SwH36v/PZX5oMLIMbuI45fkJCLFaAZR3H8QKRRYOgwRc
385Aum/d3cMTtZ41S1DbAqf3aja9UnpsHJrnssqv1poipWjL750tmia0/YtQodNX
//yDHzwO4k+K8ewAGEGp4ooXP762a+A1r9PA0BGEV/GIi2uo0CHTEi9KQUFFerxT
7ploVKkVtufDrR1OGzbKlxTMfjHDwWkCFGRH4e54naS4pjosay/2SQHC2DXpPHRp
7WtWJAMAg9BFWDtdcT2+xVxrPARcnP0mXN5XTQZr6VnCpDkXs7r+kDU3WoyPmxqp
Ew2T3zEbDkFEa7uOWCAK3boiwtkWLt+Dxmk5vv3T6B1RFB/E82FTNTJYg+PGOKi8
FzNUcOlNjxDxslZKBHdnfgkY0eyU/KJ9ZCjTaG+VPGj6BYAmn4fTTIlQT9HVA7wq
7pyiGOfc06QY2Q4z7im3fgR1jvy+TmTCsinyj3MBvICT9kxnsAY1aEuMplWPm5l7
2bytzGo+O+FWZHQDI/Yf5z9jae5KqyQyUmtgOTTexzMhSmE3coBltYD2cCeUwWWy
uwfRWDrBG1406iu6EmevTk+Jv3jhxSQ+PSm9vu3qHG+ral+NEhaIGT4kLtuHDy5e
fWyoNRI0VNmQPqM9De7i4EpF2+lbslPhrP8tAN4A1/sUgnO7Itzwm6E9TIYb1eCP
CDXMh/yWyPjZ3LZKdpGC+POmABV/qIuZpLjqjHCscqh+yf1B7OKyQwucWWawfjXg
1XxiSbkwGRwm2xDOikSK7P7n9+Et/myW9KRAUZ8JCb5iqtJNQkjoknEl84q9kCM3
TDvBFK4QVnhPsQ6C1O4C3ofHzTgEUq/qJB8+m0UuhXXT0du4Uy+mw6mPzCy/1j1G
GfnHG4o5i2uofiX5/kUn6Ci2bGpxHQUQlq+OqhTu9yRAGl57a7HgV83oJez/E/EX
86Ryd9ahxX1ajwJEZck4udvMSzCpxFTGp8XOmGYiY8slZH7PMmGhL5Nxz8lLjjnV
VZEp/Q+aUcU+5D/Lk0hecaeMIR2yO6sz2YVraG3Y5DPanA8fWu8CMqGkzLWJhX/D
Ln/NB6djRRP3QBgn8RtVZm23bPBdKEyhTPFD4LZbUkwpIBB0beTfVPsoealckPSg
5G6avTUe5p9N9l2w55DF5/v5a8ovo+hOikebPOkgq9jTGGvNBSveXAYGt3/dwrNb
7GhL5qGt2g0+OTeJDzJdJrbkHxvCAAQMHC6++g4KSOVfgxfN8nngZoQUhDe8uc3f
9E92tO7vw7q5NxGA+HkpJ5I9szDkx8vqA3dSXA+g6K94HpFkL0nj7vwva7H6Rimm
fR8n/pm4gnOotrMwCTPI4FEw6CnqLNjS3cj1ceUGJuMwrMIVhVhqBJPsrINIjlTD
1QfRMMC3w2aTGKMEULb0IdhC5Ef/t3KnaXgSsohoQbkj71NETRIzWD9PqTpgistC
M1akjObAVYMNeAxfHUNSeNVkMQagu3eCS/3w0i2ZlLQW79PYLY26KcZMiARiIfWR
m0PBacAJTTkVQDeyBoUMHdHNnl7BGSRP/pILr9NgQjWFmN+GbNxggrePkQt3y6UM
E2d5k0WG85IY3jTWWV5wtcyFJS/T1q6iiOYiW1uhvb4XCwHYXFuanDwItwoPeUWj
460TjFlTUalf4JYJUDM3uByD54nUVloVx/9bXdBeXan8LRf0EhloNmqWKlMQCUIa
qEvqEiX64aHJ1NADunF/6n7Zoz/D9EJElucisN2YcWyH41PVTEpDU3HZASXUvZvU
Ko5rjFg5bU6X3eE/MDyNHpgNO4YjMbRVbT04xFReG9rcdOC6r9JCet9uLrUE4eR0
ZpVYKgRNkPeXmedE8n6oybyaKh3VWrJONlGweAXgdNEw8/kFtG45mZYVX8b8hzQi
rJI0EG6WgbLEeUY4cJajJGowfoj5QRaBCYvkbIotO86DHl6EHI4shZXkvlr8RBOe
aLTVsVDYuzefQfDf4yAJKeFLSEvK85+cCxsxkSNh8e4jnf2hCCJ+2kBbOFv6R+Ys
FDHtLGq8dpppn7ExTTfVrmcxV7NJ5+Dmrc/zbE4rwChcEO55BeTlCGzev0GRNiSd
WhsXGLAlF4e9Re5LXy9Yl9wZsCyvkLeASY9IOaygd784JHkxBPhEn5/fzcTMHcGl
Ooz3mjP1mDM7PAQbzpHuRmGReSYbOFGDeku2UiKrrEjHTwVwqrpR3p6KNpP+kqHl
GwOFBVq2EwwkQegrqASUY5SWQ1pePh1RMoGnak6eYjgyEu3GsjBfIPsUH43tC5+m
FmFbK8J4NGblp4E6k6ULOUvabB9PD3GwQ38mi6vmc6dZVShYdr5ei5OBrid7Rbt3
GIRC+qpEJMasqf6+iTuT5Pu23PxC0ewyFHPrRdMRVS8qwbddRcT9X0OQb88sqUKb
dQAvCFrF73zLgC09fNN4qfkWMltaTnHWYpM4AdREz/J27f47aH0LntPQDmrk2WrO
JKq50mHkFWnZlzkvv1IJSHQDEmecBNidGMigwekswv6JiSa/yGbN0uC1f3KEpAS/
17XCLmYPqvPsglAOfc0ZZXkvLduJx1LcphnnGEspJhkbdJ6ncAyQ0iCQg8F+xyyt
EfvmwzOcVADGFqiiI3DQXFnh+w1T4DrsZZvSj4QEBR6RTYIdfR4G+WMOjWw6vRYI
ZOSajd5jRG8GxgVDsXl0pUT5in6ABoxFF0rTch9N4X6u51oWGcyZe2cNrkZFrEXH
af3myEniqyi+y1gwExyIoXYuXydqt+7ikIEx3Qz+sQ6I9pkxm/3g/vg0zmBCfq+T
h4xUfO9/iXF4N2JbAzely5BqsxRBREOwq6nJxAgSVfx/ak2evCtTz4ylcevyiZIm
BW3r4Zp9J25QYXZZrwTHfKP+o8pV+gSirlB/yXjPI9dH29gq3bAEimlmUTlbY33r
qa5VpM72AWt1sDZrss15CUh5fpviTOtTXyS2kkAQaz1oU2nCaI074EmArvbPUKeq
WhJGb9MDZD9a2wUsbF2gt8RJpFUwuA/6pTr6NwIJfp0XiyH3zfRqMLGoEz96XyWI
v5QDXwESbNtWd0UvkaZII5naCyyhxziYlsB9XVicRhk/ICmiTMjkl2H3Hf3dPW5s
Vx0+NfYeO3EW9T5IH/rfshrg6wCzBiyyRklE5PWlJVTXBd8yi2t5h6tFk07/NqJJ
vDAEmQOh5V+ZWIkkS8yKC1pSRLn9/S41iz1KL0LUkrXQ3RHlgq5qoIocyZjiHrnO
zhynW37i8DrIUjyHdH1xil88t6dLB6GSzyWXfeQp2oUGoRtqBnfqHCP4m8rwC1Ov
UYqkALnylQyAFUXfzhrlTWxCky+T5uw0nfYpLh5ywcYDy/NGuhUU7EuFfEgg3iPE
9nyKrRliQ4zpZAhVwgy1aWAU9FXJuBgPhn9R/fyTEA9YZ9SEW0Aq3pfMZwX504VF
IWj/IK6pmlUMohLzlxgkzPGxsuRtmXEhE30xKAkG+33hg0fW9FQoSzsOOZW6py7r
44X6mxy+PjSo2z2RVWVP1qmRbt0V2GzEhl5O/K5QTA31IzE5rc63i/IxAkyN2aCx
HqFi0ru0ukz+wx6l+XknlmOzbr09ODLXWGIDwzL0NXSbqrQvNmYQpaW6Wq9BqpOl
v5DdDArDJfPIlAtOeRhY9A7PTHbJp3N3CxQb7PpwmmsWZkBsH1kKg7VEQtSwOLWf
Ql17Xj0HsSK4J5VneoCo4we6YXP0+pNKGSm2HoaWqggOhfOUZPmxN/qgZkPbGjM+
ESD/RIRKSzITA/nhzGLz08npuWOQgcY7Brqvmt1rW8ro+qGzJJfaJJNa+uG7/WuR
dvI3YSx6wPxFLcaqfzI0NhPpEaKgK+/bmqrxEsFJb18DJFsW4jpygzdCdql8Jh+5
Tb8rdKX3XgMNy25c7l7pgiNQ4JCi+HQcAW6rJKipO1oG9DMk6ZKp8zHNb1ICay2x
CP4x+6Kx54OmiNbZLe/TSiTqO31fxmqwchYaCt6O8hfmprkIKE7EkgR2WnDE2SeT
Q6wwwmFkHGseS19+lCKozDWv9BWADD4ZsFaH19w1vs0ACOKLv8vdak8u/HtO/hJn
S/MADJpE8N+pQmLeEv15faKBK5/tMGIZJVKW3Oq4l8K2NdsHpjq0OT8IWbHQ0oOJ
yKJoXZlADztIT+FW3xsJemNNDVlKp49Bvt9C/jR/YtPuQTOlkWLfsFflYjwdsFoO
LS9QA04G9Or0FXLVN9XSEtuTBmpicfm0USboXZ01LBv/Ul+sWP3gk4lLH9uQtCWd
`pragma protect end_protected
