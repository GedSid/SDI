// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:35 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hiwRp08HKCH9yZHeNsi3ywhXw4Y0hY6fC8oqwsGWJBIDNkxGdnB+Ev2enlJnDnMW
A9wmVApLYjWWb5qzJPTaeDbu8U0VdydScltkNXxdg9HQdXf+mDEBanIPhQuj+nQn
E+ahbtq+/bxlHdoy1J8K/ChVYam/CTJqDZLE4cdbq/U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22384)
mn2cJamQMq319pJI2usPiuOVe4dm8uM0SaYN2klM62OeD66i7xXkfQXSL+nk5uCE
zI/dWxZRbkovookdCs85skzW23Ymn9v9hdOwx27XXdAJdsu+NtCMNLIfpftlkMGp
4ZwW57nRF97yly0E9HWoIujO8Aobg6heB7UsW6JptrhQM1bODm0m0OcombB5XL/J
q4Wzj3t9kOWfp2W2V2gFK/1AZf7/qgeYq4477xcartEMvAFuje1DoY9V8IuBN4uW
wbkE72yAS2lj1D0e/4IuCodDgLIf9N/9KA7fiGW88rTUHNnVmJEiD/M8ksZNiT9a
AmsCjaIyiafq0e3cAIaGenaJJBIKen0vn8jr6GBqVI6KgAkqBLSLvpMnwjwq3aaL
2AmyeB4kHN0eapQ8v3nwW1VSk7EgnM7mLp2w/EN2NNOTSEasu7v4jQDf4OjG+FVY
XUDTPxTPsuDHfFLdB7LewsJ5Tse2748WvUZaEydnfHswN9kQEusH82D//qog17xz
EM8zvtbJBzw0AEd25T5RlZdldudxsJgbHtmQWIPI+30kt6wKQOikZJ7UjAs6+plU
GJBR9eCP/6o1aCeDSqBIhkZAYUSYiMrfIW4dpZXkoGCLuCzrjKsgXFb9HP9PHBFy
ZxAq1K/QjRm7biNpID0qa/RxaoDOg8HV/Y5cQu9FTcyjb/thMkPJ77hOALpuX/dA
28uFSuMTOAvI5qpvsZ2pT50qdy3au7qKqoPLQRLGS+rZ6GG5gHLfo4NmmOpqq/o/
k7NTWlAuwsHCHAc1lnHZhvfc/5iY3cKfBxJZiGu7nf944OHOzcl99YS8iWvj7BeB
VABrUBQyO9SWW7aWqGLI1pOB2xstmvLZaceQ6CaQe7a0Jw5D/BR8FG2B+vCm9TPW
ZJs1Inc2y5mr1R/9qUIlAvO8VlXo7uedhbi+JPU6Y2tpxBKZ+zGFyL4VvR1yO1H0
+ZSoir3WnSfDtUvZLAFZqktHgWqYn5w3WWvYyiOBZ9gfcNvv8VP0wMBOPNPNqUVH
hPYmFgf5QmsgaBw2yhIdQGDLEzGsXFsvQG9TBpT6gXv5l6KGdCh12gOshaCHukyR
Rf4YUtuZVBMBFgy2w3r/7P01gHQQdozUJLA/afjAJ55IEuqIKVXSI9VDlV+Q0dhk
VRXUbFP6LNYVfC4SRqDDeNDW2tNMzYCW/DEpsMyq67U1WHi1/HGdfWiXHVdWhuHE
Qa6seQERBCxswqWanRjTrjQccn4213j/5xoi81vhf+mSgMrmBzJEge49azhiRU1+
0vtPcxIdxxNM+q4fEozSyHv9fEOnefnZr4ygl15MXKIw8x8cxyiYlz5fOhmvuCQp
eU452qXpvK4vs+yVkyRhTXoX4M/V97bRfsbpJOrjlUHBhpVeI8ZbTp6RKWHOd0Dm
woyhjmJqh4f2eLaVfDjzpjVV/4ws25/iUiwaAty9+TLO5Fr988Orwle1Ak7DVsil
iaTbbvVYm8ybori4PA3wDOT7rc9+S6EeSiHaeKD2Ns1ccpdgOvPO8Fcl2FhsPB3c
ygQhXO3KWSwPXwUW67NKTQWLDkruST++eySYblXUfBdGOOWTeSA8zS4D2ZjVEIt7
f7dYuiUgYyR+BSoeEco/OkS/ttE4ZoWm21O6mWXGekbzm1tKde8VKp2z5DsjMNLV
UWTrW4YI6DonMjNynjEGrs5yRrC5+0xh70lOZScMp2c1NG8qkUJVr7bl4z67Dnyi
PjjlVXleZZ+vGhcLHqgtM8XhTNkGIC0vFHf4Nm73f9tYhmOZ1r5gJ9g66Y2WmiID
hAYW9cpNKeLY9d4xnLN11OdPnzFeCvCuaaBAytmWq/UnduGwHguen+6xxRiCArkW
xFyuCoBySgb5n8kgE7wslGX35Y95WcetG3oih0EOVzIUmbzsA3RBFHIM7JVe/Nxt
Z3TceF1egkGe3rNjGEiFhJDWa52v8Gvlijalm/DD+c58CfaiczCFeaV27U0x0nLI
VXsRviHIc3TLkfcS7H/TYLnjSuU7RLW8d6obGTytgiksQV/0wCil89DU8KKV2V1l
HnDzuDHidf1qaS89wvRykJMp4GTEV7HRg/E8d1p8mrf7wl9oMqxieEmN9ZMmxEA1
UdMSDvkUdupVcxDRmTpr2q3YCxTjBjongYM/287F1Rhpk0HS6LWn24+z8xkeFYhz
x+hOpQW4wqCFN0Ni05LMygSxXJ35upEtiu0f0cutJoyIQ+HYtnCWKR5cqFaMB6Mj
MCJ4OWDpnx7FdY4mCaRWJExDSsyRX7CBk0tlCgRjH0rqAqtzMJt8882EXfn0741b
pKMgy3cYvvDY6mY6xhPgt+aqhmpltR93gssr/zbH8D4wj3Uv4WBlMDo3D8aUx5gd
o+s1bV/fJBfAy62iwCQPVKgDdWkRR+WrqWU/mkwQirdZ2HnouVnBKYh+sRDkg2Dk
4TUzno8mE2FHTQ1ps+keQJEfg9rLikjqHDo0Yv5evRur5bANHpw4oRwTNDzUycu7
3+ac4Tf30Roek6fdncrkFlq8OLoh7jmKbuXwO6laIN2yo66reXt1vFDMK8j/OpFD
1tPO/TZm0w7aDsum6KFdlqrXfBmCkODwX8T+EdkV7OUpLBbuM1UjhfPlSX1I35yH
TnjvSIQ5wUh+exTYcOCRrRs+8h7yguQdffzF4Y+StN40GbTWg6s/zVET+pGctf0j
hYQHgSm8P1WjGIqn3a/uJU87VMMvRbSxEPAyi9egatg0SJOMLZF6pk8o+Onnayx/
zKNlgKBKDAv1voeug7TGINA5d8pkA+u2iH53P7KvrxlYqte4K923krQj/N04VMMU
NDXSN2ZdUP0CjggpDVgk/fK9ThODqUUFnmuIaYSbMtrCkPShBrQHZQnHHD6eWa3f
rjEoJqteV0KNjxdixE70Anc80xQj9Yon75H3y594olqT3c0Kj6W1OLc/CYjawQAG
y5AW1V0CbsiXHFDVhTcFnzII2csCs8cjCob2xInpg+ZeufoSRdVm7shWuidQbF5l
tnbcQFf9puhE8sFOzjtLzQ/cjLuE+7MXNxjy1GmDkSnjb+A/yFkCbaCbm9r2bNng
lJv1XDiI+ZoOokMQxvusewrnkGOsGURHEb0pR9dKRwmPDhUeVCvniw6CyqjU6jYU
IZQCptPKMmOCxg1L2bc1Nz/ETFP9SUVUjpYmlaC6a8c8pttBaJDDLC+4drQnl6HR
2AocHhIRT5MeIaETLosXiG7zPw8rGbhAsvxC3Qlqvy6+pFs+mOdBhQ/ruISoKAwY
gLLiF2GLKDzdIlVs+eXvKxvSz5nWfq3FnEXo1SV9MYgeL6LAVxvJkRh1HAanAndF
prSCRh2blfnjokEt41AXxLw4Bx9Sr7l5/cxPAOGGqyTOJ13taXDyWJiY4OWSd7Vq
HOiGseWRfnCenV+cxXL4UdOFLdRJrjRYBPRz2qCU3WXibFnm1H4dc8X2L1n6iuFY
6BpvjrDxNbpOp+vfoY/NxMn3BTqY0hgmq7VsYtw433Lrb0BZONq3VjrbR3hmpHbC
UuEV+f/ferSPDyYLLhahpUjd2k20ldDVHpZUWBLImjNeBAtPmWCr/yyY0+ZYlkZR
2v/k7G16H453fVxpAoZHgZgfX3D1p24fpg36wY3qgx+zuB9OhLql1R+96SpmVyIX
hxTf/7Inf3Z6SlFBXNkxmKJP3FkCRb78/ddcedXMwAJP+Sl+IUrc81zjDU1IaAyJ
TChU6H5tmJRvyt7RzEqtIoHmIAt5nlRpfwtzz4i7H8NQiMftyMrycDsPDJwwxe4C
JmFQnraGoxRaAmi6d32v92pfy8vuLGZKD3907N+im7O4aHocLXbM10PsVttBg7cc
/u/EiCmj8jVZhd4QrLmfeoQOKXO+z01nI25t6Wt04goV5pkJWWjrrlqVXkJzqnJF
/BTrVJE/YyDLIhXmsr1mZ6eT5Efbhp/BKk+s1mPLk6IVOzM1+9EnstEhOfPKDRP5
p3g4yi+9Cyy6mw39PkoKiGZFeU35b6drxT8K1CFRqAIXZQpA9k8kBFByM5l4lmx1
2gbEnha9qqUjhbg08lf/1rPJqEmMiQDnDkz1RJ7mxkuHya2YeMFy09hW285+gjSj
rjZQGOKsVXanS8FBR/dBJ5ZdTtSHfdNSHo41YgAYr0E/NMCTWKJsoVlOEIf+At6n
hReW1yTuBstnAgGocifSIlpNmtaTJpTe2mXV68BfBDZfwFzuBreTPO+ri5bneBME
kEUOy3RVXt1KgbXytuJGLOQ+BtrAAeKbK7fiUlw4q3O1rqhRtb8/Y+/FkLncZ0Qc
JT5laSTQWFgFeFQx8yICI3c9hkkHJO2iYMP/bRRFJL9kKpNpjVm4NB2tlQIgSXWE
xysWaYl616O3MlaLiQB78ktNeFNqF44Km8YiDFyu2EYRZ+RV8xKIlaIjFaHFTLV6
pnsKiU0t5JH/9++djZsabyjqIj4AB8XOANsNRaX3dFCRK385qYaChuwnXvGU6GxH
j6sIjlVYOcqr6J/hw7IfzNAtCg5ykqvwpLrT4Mskkbqf1v7DSyKeEqfSHyD+zaqk
tIyqC9YTT5qMLZwdr+6PLY91EoTf8+CkMPvObp9R4D6YSD5fDo06DaB+lVRX4VUi
PvIhj+I05L/rdq5Y3jMDGA2OPHooA3IXspY5kiyW0VjPOurpr0XimDmFzLylIq1l
AXSad7o4BB4A42rnTT9SpIEfjWN+UvoEHtYVND258kpN9ebRs6bFemOl5vztxm3H
WSmsoF58FSXsP1HhxeMeJdg9C+43ujimDxrqA+qm7qkBGfISjONm7JbFvhTEAGyc
OCYGCn/3njCDOYlagxQ/y8b0OTglTgenCgSliVf4jRYlJH8eCrjaiYd7XoNSyn/O
NixeS8OJCQzNNAbUkwLDBtbvKSjDtZME+zQUOJqEMkEkY+2ic+WMVWTWiUZfSuBu
SO55BxwBdhVNVvFWKecTkw1U6zP4HKXr4+DeYSnbE8KFUk6sJfI+JFpDcdbT38HF
0jkO9ikmTyOmnNBTnk1I+tWhKyvRb8LiX0kC9dAYH3E9GepppM21T5qstq6AiHq4
wSeKeRp80KZfIbGIGSj7ymzmBFfQgSJeEZdynyUBtR6/dQ0mmCj4VceBeqQmOl14
HT/9GMsnejnWx97CzVySqtuV1YC7s0JEEGcUVlqTo9TjN+Zu8BLMoJzfOTWsI13/
3h8pVb612mKYuINPnNzsrPXvQzomrqlcqtu3sMmwmWAXxy7M3x1KufFmWa1rXPRH
QILd+lv/oFhkjSlsK/c17u7xId7V7v9DU7T5BkLWtBWoS5PTN68ei+Wc/odFWRv6
yBawjCLP9NL/fVukXfR0uUiTm/armSt69rMd/CWMHK8MaPzxwswO3axnaNV7RJT2
6pux1qMLzE+F6XsiQOzUrX3BivVWgL99VTXs5SfxbMgtZCPamZ1iheIqdBPXu8pe
z6lJlr7L5yN4Z9S9J0Lic7Y7EdNhS8ySgAYGxw+bVOevfEWLvj+qidqeb06CzIHs
M2ufvaAq0qqawYQaF+0Cv5Uk1dAwjlsgbxXA4xLfecQ6x4nB2dxIJyxMQbtCuneO
v0neN0RXoEkxv/dodJOHWuDhrsRm++x9rvBn5hHGseu5PeDTek/wq5Ry4rwxWqUr
lmhDfsH9IyulNY7GGC3+VQu4W6AGNYemexiHfXFXDzxRm7ZsVh+07amFgltkQc6r
egbeLZ30XzrHdrdWUvkJwvnnTlyFlU0fYYKGmuSJG6grbky6OwoVLQzirBDjf7v5
FFCxcpJUzY/fXahp78UjhCSiVcD0kjorWuasyGZMxI3G+K2BxbNGMiwbA64FS0L2
P4UT5WiIUjzk/XabWbCzxht4CdyFoQM6kq7cAW6oDj6jjhhFE53jP61CKej0clyg
D06FCbIUbJGi+DXUe7ca7+LtgR1K0N7l4+vpQaThrRsrCHHDXvYpyuyyjtt5D/YQ
6aEuSiHJ+Wwu0FNZBp/i7L6nmjMXEwpKkJ1K2VpcpS72YdI3ptSzmjGNrtMETBqG
SgeoDmXyGCvd1tcW30Y8IJ2jl9qUcxzazbTi+l17Bo6mT5pS0GKoU15MrbAmG2vM
Dn9ddwPBUZ0rjiab8KTF+RQ98v5T6byDGg152kBMhI+tGw7r4qMORUtSvi3/HYpD
8Zqygr/pb1/9D17WNtrE33gMSGSSNU5WwA9VEmSR2KM1Uyf9TFTuMygkFgI4ZsjJ
g5LsuQM6bRBZFbJSI6DBtfvqtXkbt6ECTZAJs3o9ewo3TN8GS8fUIVL5Fd2o560/
YvYDqcYbBrnywTVxdyU6EbND9rPievYl0YycPxZJSzEiym2NoRHJ4NCWAsNMLsTa
jZxEcU/oH0PEj5d/uDKaOHAlztCf0IfmjQZDkAp56qnhlznHKFMTC6VU01u29KhG
/wDk0YVBw3JAr7Qwz/kSGFthdf5zg2MfS7EZoA/CsD6wtAbTRHW3pL+VO5YGht6d
V7cwwWiOvPo0BVlfVKZnF/qbS+WEsG22uYnJgTETQWgOynyspqYrLLRhRNUyTZVP
xia31bpiv6sym58GIz5wfy3+rjxuLEhVTG17UK33MhJR4vQ9ad/dBnvddAO7NjSv
RlcJjPOCj6SvJON2ZTOean57J3vFZ16OkaaImhmDNCpwgdQ2ltSrEyCx7pZ5Z7us
eC+axSojP1xJzRMlYRCL/ALEVPkTQ2dn4LGR/cPbR8HunkRL4x5XOA7mKMZZJpyz
tv5VMk5tUVrvcgMQiT6Ns95ARgzgP6G3Myzgf4/szpgi/sHOpEP+h4zEl0hNEl5q
9KiV/lh2SXcEiZnAVvgRxP5DEdoEZaDqZRFoxyS0n5+nYG9OmGm/sBlFfEvplmYg
XCchIN1syexhywZUUZjmwsxPdyHIMVcX6TCwyFldzo7pc9szWHTVG1x/i1Ve0TMb
m2MJhE9Gfq1JiHnqUR7X0AJnzyvAAKOnUZSTeXrYlydNgmllrrZsuDJs/XxO12HQ
I2Am+IIQDttp5TsqlMrJA83sb4tivr4aFYdSQ4HChc1cK97e7tCK4GUoEj+s52nh
59MV4K98QveDZ2hnxRwVJor7C/wPbc1CbcJypk26ntqG5Mhe/h8DeoKAnB6e3a2V
jdBBUSvolZCNSwnSacH1syaiqQr4+iudLXJ+K0WfjmsUqne8PBxSS+8co0gjftTs
u3iKbtp3zsGrt7JxRC6m1yk/dnqzcIm+4GuvizsSpTIem/vFAJ/50KhU1cpPZNu8
lmFIqIWnA0jUoNiWB7wQBYBWW5m+Rr05bvyb9HoYXnA09gwb7TWWnWWRwAaKT74T
1H9qxCFAMscTAg1knd6pQilv040+O4N3IVmxmKfKnWyaWYbdE0JPMQn9J3/TyLag
g5X+J2ClOyALjT0r8AEiW4mrEAwHxTltyDEzHLT+6MrfKdicF8iKKYXi5t9hhvh9
9daewdPc4JWeqyKWir++t67II1snuUSECOhM9ZhmZkQwVXn8iFRUFIiCqLuyCJS4
p+7kcI2C60X73O+2G8KddchDlPvpwqIi06eyetE6PbJF3pVRWBBbcTyjVaesJJLg
1R+oF7log2JoeXRxrWTbG+gHghcJvtSa5aLtNZrahekM3JWwD5fAM5vBm3gGNaXU
Ywsz2AIvedkBnHY0/SXxEpO4TJImgW9dNiFgZkrirp93QCEugYIRQgjGjLZtPxAT
lbRuLwBEo4VJ6U0sv50FrGB2icP0im7WgowHJg9fHS3I84MSXcIatK/Qv7LkO54y
NL1ZrSn72ENsvdg9e/R0Wg/faaDozVC/QGlZVb2NAx/d4GGqxL7XSrspekzA3IRA
loAZpXe8OsPFeI2t+5H9AVQOqv6PdPwyaqKBuxtV7QZTFHOQ+DIJOY1Jx0QwguJU
6fpM28ZlJko6ymahxnCU7W4ApWo6n3eD+0OT+3DUFb935dzfoEgof6Kt6rRrpgrT
3euiAfpG58wawb7NXsIuzKTBsblHGjrS7lLlZg/NPiLDHpo8IF7xBvt5PKF3rpSY
944JsiRVki3PuD5jztZbNiC/+zoNoLmDPD1LU88iHygm1prGw7bwg/7yDEZF/7nf
eWPQ1fTezzf/e4MzB+vECEEf9Oc/OSGtOjbXO9b34bS6ibzE+JTqfjWnq05rv5IN
hQ6i80DJhBRH8uE2UXblgb/bbXDTT0LAxXNnFA/N2jXuogkAkRliC7KlHFUVM9/S
+wQmwJ9Rtp0QAQOwvqS+NBn274Qm2bn7RpI1N6hNbeY+/w4QgfpDp9eYdSxaF2n8
V3KPzB5sbfYGuZSU44YWjRUN/m3NoeW2zHcQdJqfhqbwpznhwMqZtJSXNqGkPjIs
G8htxB3mnpUHrwJM6KuKHUvvl1m27J4DyaPJDhFwZplXwmvsiWlF4yISvkX2tx1D
ggcVmqYOJSsqdDFeA1AiP+GNEDf3b9JUAKjyHY0+Ub40bFClnxiteTVTW3adCFZC
d3eWxbZ9PrhQE4QQf7KeC9wXu8KN/SC5ShmzrZ3sjQCgt+af9KK1KaAbRV7+9dtp
oaxe+FeEXPobeK7VdxKymSPXSBgo/dlR43iaUe15DafuxH1m0IKhk/C/sSK0N5Pl
Zns0/l4ADtm0f53ZtA13Tbt68z++tV4IMw1rkZvBMYCP38nnE8N4vQND4I3gC+3x
wm5hIWp0Nw/+4aH2ZbKP6IlaauesyxelKO5hPHJoyDsGqO3WmFtM9nyEOBWYyCjJ
dEGnxwhuVpwHbhexaTsFA+fat+L4BbjMRlBfXEFOJDN2EdjS+844rmaQg2qif44S
fLC8qKLWEMXpp2WBYHcp97duCX+mJTPLodnuXs3DwZktAJLc9g+vNsL90usC/QnB
3jnJXY44R5oCPLjir+LydWRDcP2MEvgFDoJ/JL5R5hYUlbeJYQdcX9mOofDD0FEM
VnPshlYU0TdjjbWDOpUsmqrLzKB7KkwCovzZrDMMpxA8EpsZW9wuBSAoXvdmzKHF
isD5SdzZwZBxuah9N3zOZElfBSfYCHuMQkSrmS4XYbyprW88kPflMD0Z0oppb6w1
ybeM5LRsDb/URLMAjmZvP632tHyIdEpgk0M9YBpK1BYlNqQNJU+zz7C895XWlskU
6y41XMY5mNfKQGoPwnEGYqvUZW0yntfwK2/LoW3vm3IxtIgn0TiqQIPxUCv44IQf
QJiiNXMMI1dvXdDx2y3MKcq/RIx+deWrIVllZ1dkd7coGkHvYxdhQlltndYgu92g
7o8SF/Sd4QD+CwuaVKNPbL8lv4Zuvhj3+PMUSB0cVsI+gYPEwbBrcNnenKMRIbzO
ixpkrSs8IEyuY+uiaLZNwjOUZ0feB7xgQ5Q4m/wCTeh4J/li9z2+GEVpOqeoumHV
OGpjdwCshP98y2lXbsA0S2hIqDNJdURqJC3nLLUp2CGa3mL+RDWIxLRJ4WdSbdst
6qJype6C+oVEZlNbstZKEx4aPTAwPAM9U3eGMVKQXo6Lv7eErnEqF4iQHwjG4MC4
RRpRQneoyVGfOn4TZzo200qFnHHLOkfyOMBju2Pof+2BrMBnRlYX4KnLMORPfa7Z
m9y+D2uMw5sXeq/lFPScz8j9AyBYvFALWYFGqcJnLo1QGJ9C+7lhnR+iBvdjkY6+
avumZDl7yUHF6iZu+5rQrMx4pcjacQJ45R7btcI+esOwL7lSa4PuB9Rd0DjScR2Q
PpKMoVGR0w0/i4B0woi0qEvP7ruZtOOzRcxlsK6bpdDJREDsrbVKdgfhmArbq1ug
c3aDx4Iq9Va9rbcEPSH9dIhUgF7f9FPvcaE/6wqgVLUo0gBtSxDxLRKtHb83ZMFP
C0JLFOcrTCNK38RAeNoasbUMOu+EOWbQ9AqZhXYX74KiDTnTQJ+GOR8YtFAzRYPC
H8LfAv3upl+lY1C1iX8YTLzzEHeqzjiNEMxlZ/uFHx8Z5hWZ+rSew4+vngek3Y2b
nV2ZbTGIBvNk7TvaRlVZV+Vmlh0kjJnjlN+Ux80RqilYDiNUNa2omSn0FcCkthBs
TtTEuFJpZwaDvhwR1whKXAL3X3cnoWIhCyT9MJdrLDBviSa+/PXH8Y1zzZ+yOyyk
y5mHRCUk4yIrwAy9oys4JO00JPvJ6AAK5EzrmVrioG1lG4/R82uPke/2B7TBU7Qc
5n+gVEhOdltKrvBeUo1h2iJVK++ZAbiJ2h89la3KzLI3regFO81XWbPr5IJN1Yzl
LjlD1ehLMVaVdRv8V/9w5kxQn9ZbNWBWoSlCSQAZqfHm1R2rP26LYn8ka4vyhVmF
953aikjWptyuxfrpjxvV0VJelZFByE2f4d13CPZBEkBfkn9mu30azwN7dCdMpgMq
hv7iocPPyyK5C+3AdiHMqOK5TTOu7QdajTLMcdB5JtjWm6oXSLm8OtNllqTjeixH
uTbX7ZZ1GK1Z/JVZvPEWnY9VFQxjUV+l4SQLIUINVBTAhOq50vv3ZdEeTBbIgGde
tYNJm7DE9NSRO1hP4VPUkETBcGn9owFkioDrO6DwtdVM/vowr0Jb5wAkVrt0YEwt
zFKF+0M/uf4y7lbRNwLMrHG+kN0TP2dQkx2iOPPr744xbfYqZIVMRb0ciKBcGQoN
SehFw/KdlulOqu31Cx7hdBEELqx0ccW1woBA2xY8K8qBj49JqIFJNfjBKjJZFHby
uT4KzVKoKP3MJ37SlRQImOiLodLsqOnzko5wWDfYh5/oDtgmBnW/bUFit02BNl9p
uqcqEeSFPjBtCV6djHRusBrnxAxGv260nFXIB9H+hIkOIW2PIY5zZz+gWhSR4bW+
128DvVjWU05e1OeVB2s5K9ziRKTu1Twl3z8FlUqI+nspok0zlbv5GGfgJRXk2STs
dEc4F+Ubb4HJCN8mzKIOwhPcFOqajlfHFmLrriM3Bt5heBm3ACmNMgsLyl7LMiXs
S9RRQmE327DgKaJGevKic1IxXk0VAb5pJ8FMEyvtpblNbSdZ70nKRKVuc49/2jZc
6orbpf4gmeg3wNfCBSMHVfTmju/t64rfPfn47hukJx59n2KC5MPtuaRhpsp4YuDC
SoonoegUNjq8W9rYqlyxAr+mRa7wlc+wLe5fcd5fMykWfsxmbCLOtRwYZoGaA63O
X9WUCJEwHbq9c5euB/46F1SiuK0bokQhTxufbQ5R4xWBZmcd1zquKN0+FXj9yspZ
mWvjUyhj+rc4NSiyicxe5J2FUSm6154R8y7EWTcdS6zHuwvKOFFg6fyBbHtipUWp
L/K2q92Ic+s10QLBWjKb7eGb/bgBK6IisCw8aUP3UWv7Z62PKro3uRjjbchVGJQp
QvfDGzjCCjybvcPBfpOOd4+mgOiZdehfCV9/BTTr9ZYZd8wELAEEfdavu5k5nk+4
iul6Z4Me4lc+BTdLQDjBtvpBIwbrIysNoq84t5YvjmsGuu09V/ZELXW0U8niXTP/
GdctDc9SZHAXOu5jDuyyKtiiVzg0YBHYRACHnpv4my0bnpVkWV65jS4LmZa4CITp
kuM2D3kOmKFwm0kG5KNI/X6a88VqxR8TMLXCI2UPMBNBpmjfPqCefXRR2cDTH/5O
aV1iHlCWss9DtGIus/yae7ub5RbTzQp+mrh0NIrVRNAOIpsY8h0uf2HNujP4XL+U
18E5kkptzDDs84h5AhoNY0YP9azxP4C3fKa92AlYMbUuLcySYeD6f8EHJNtifnCm
8XT6HOhEE7QG5uFWV63zDhT4nxW8iPQvSe/KqRlh7qZ0f0xDJwBfrdSsFRs1V0Qb
8x1glfJYOS5wViyjJUB77JQwIghsNJo95QKSPnN6TYLiPB8FJGCoZaOocfCrRYS+
U+4pMpxZUnVre95jlhRcHXWQNeqkPswBg8TizPF1NJX0Kso3jxAPMBtkXfEUKRnO
ZXYDvqsEC+aB5GONGRMnQp8XDOwk5CsEH9gdXIBGU8XJdM3SA8nD7Q/ap/EIK+VU
09+pPhL47O9HU7EX8eeNGsu/Ddl0E+Fl4NtTi3iGSCW/5h489lNaOmX5vG4vPgpD
2eL9O2+nKb6Owv4JCfVZtL3xRAPbXvIFHxBEsizdgQzX8j0L5SnUr6OlAtj1kLqV
SlCLQhFKonm4thvCK37gHf8XP9K3m6cLiGi0+DRX1PTIS7gYN8AA4Jj6eUEm1KiS
V0vLfwSIaSxbB9GPScuM42If+hjG3MTRC0QLL+lEl9x4gCdfV8RA6fJQSw9xCMXC
Hcud0Ae6KnQU6QR2ITZ+Wg6P07FBaKDzi31TTQmn6R4743lkfPvsvDl94vu/Lb6P
54W+K/15k7vjLGDCRzvVZBHqYh9vFBsWjMNy/vUhdlYSE2kC17RdAUZp29cOj4Sw
CtABME+saAY+TJL9MdPfIKKB0q8W4Leja8WKlVqEj5LPfENHFnsTJevuw2hQXTWh
30KotN9CeqAu2dgWw7Hq06QpR/5RopfT02pY8CYAXFXVs1drqogzgdiZ2Th7IdCk
VwGLOEAWpElTJOpROKrlQCBXCsRN76g8ssYMUK1OPn8smanTrpOeze0K23w29Lmy
M3F3UqzEYbwuWew5qzrqMGxt2tXG4kwTbgbAwdHr8/emiDk6bJoQdKZfyc8n3p4a
hrKgQRq1t6uPo15j7UAXRlit6aiLgt/cgbUhqwi7UvQoa4pjDoQAZh1NcIqiPBqc
X9PuYXyheS6SRecEUCkdum1PlShxoSR1Rb/boSIGcBHFUeYm1viWfgeZBbS41b4w
AT/QVjHIzugsWWEy+E7ZCvVU+4vx1LMO+b1Gk2HmYq/4CtgB0X/c2nrdDXYvStV8
ndEK7h32cewHWW1z6Uvh4l+xvQQ9PLLr2KTaAKfcUEpno+fr3hAYa4a2gZ8y78Rc
tL3RVKElkrdR9iU4qbvRdmI0Fv0wKBaeR4+3CuoLsr3SkWOT73qy3S7Pm5Q8/POi
l4iysmBRZtEqklqIci81bfHF+46txROGwNn7w8OW25BQKR1BRW5/+f0FbnnTp4sm
cLsT1ky44oqJjv64wZam8APLT/TzT5uOQuKHD2C7siT2ZHYyzSoTEIF2dACS79N1
5ocLIoTilatbAGQITV0cSjvI8D/9vGk9CSBFvCvyHsSTZD8oRglbK0TQ3hojV01E
bcun52XX6ei4I1beMep6uF3DJwtFKKnXXwdTNtn6u6ifT1eIVsavjJfOefOhnRAS
+adbitCGig4pNIglSm72q1OpuzRw9G68zJ1Qlmge46OB6txAdp/OQm6nwIqBtP/+
dqNKZNc/7CCnsCqrSd4mH/mhKhqkZ5iLKxL3Eub/1AJNI0SFpnP9DP0DsXkqy+Ld
xGgcKU1hdpyVsxfZHYGQahzxFpfu+GqJ4X61qs7wg1vjFVDM43VY1OYcHexa+861
WxmcX1c01DGvOmANoWMHlxd4Gfi3Ir1opZjEDbf1MTvLC4SLhTgLTtcZsVUB7FgY
qy6LcqUelFcc6UYeMgAgPPJMMY+olJlMgui4PuAVWNzZa/2s0FSNxqIjLczPPJmk
2kJMVgrN8mAXDFZXHeG0kHBo4KpigZXwfELVVQ2ppffOXqKwrrawAeIdweqRDmMw
dwb492catBPDF/wSW3d2ybLbwd0vnZcrQWUG1IikaLmkCocUDtmnkVnGn6NgAQvJ
MRXuKNKuJfD+FdTM4RHKMm+Mqt6NosYHPgw2xwWwUaDtces0/eR0TnGlQlKIbJLQ
CBBWkkBEXAQ9bFWOLlx21T819jBWlNrkDba2zJI8nyvZZGgfCqPE2n65JuB29jd4
ihBK6HxBkE8l0HsIPDy1IeQqC8k/ugGjM+Izg0TvSO9tqZi8ih8iUE62PBS/zN9Z
A5NJjnQY/wlQ8MvcADkPCgBMFrF2AIU2rutg87oCe/0zmoPs4el2bG1dkT3MUJZi
w5IHzfObLOKhbZ635wGTrgVs0ptd+sf3QDZXJ36e8bjk2IQRcLLJXQMQrylkJZ9j
GMIE3yIazAGh8+eZK3uAqQzqsr9WrczPslEvPdCnh3NIaXNl+FlTjF1YpwCrlMhv
B/KK2AgEqGsQSxiV6xOCrIHCy2W6J+foxibWUNRGoec98zahUcPMPY3ASsbauoq5
bjs59hUqsUft0SL9cEg7yuJTdoNQ+HQJPHaDvybvjCaEzRUIrxEiK19SGrsnPUzi
XVuL8FeHW69d5Otf36FydJUryT5b6HQE647+Kh6v7oEw0z95N2vZ/iWo6fwQ29/N
WHVYG18k3XYKp+2GVK45nyVDIAFlImvKYiF4HVu9CRP6aoDrtEj5dQyHYNGbC0VO
dW2p2BbRVHEWyDsifpCt4bQL9Rq4Oygv3qo75vw9NDW/quz0mnguS9lCBYvVYVe1
ZKCPuoGE92CJCyr6LNxBc0d2v2NXdYRpow7rFJ5tHLEhCZ8Bpvjp9uQou1XwUAvK
EyoKFKNy0WdOMsM9h+Km6nnnAFrzHCxBnXDmOsm9WAbU6WhJGTCrA31i2tF0QkGN
h5Tb106BoYKkZ0sDex5Jj5GVxYECc0qpiXG+bJMwyFuzpSiQRyws7HiEQ4cqnQWC
rgsORoLl8EsSZCLuw4i1SPzOa7367dUZwKflSAlEIWWgmevxnvnFwZ7QYnrAkTW6
7gK+udfNEaWu8w2EL1UmF2wFMRXlGtshFGvo1EGYErNrngv8hBl9ok6xl/i2y97/
9YSl4lCBrka3AWDuG3qhtiVESS0R95BmioIbAls0KmVWK4+xP7VD+TC998/pa02z
F+nORrGeOLmzvuK4aYi1/OlkuQ3yFtR8I5nI27YLxPglfBfcBH98h6Nrx1HoS7zN
pf+IVF9ZExrLEn50UTF6wfi+P9/55TvSTmPPY3nWs67kChWzMwoQWwrWPaoEVHYA
3yPd4jQMuzLs93TD7RhQZDi2Owwkp5fP4RgbzN4Qd/FJZQsmZsqp3+Rd5PDMvxzJ
uGJzR1lEyZPa0Ie9vc2uVMzFV/S7qeQD3Ooq6vG0SbpOD3Kb5p5T9rGuK2RTYanZ
l+8DRoFCBMw8HXINu+2aP0IMn/ycSoOXsaHXkAlgvWpjIuxgGdLYNUYV8LqaiZee
+/1CFZHhfNEVbwVhryzK0cdKzyyBzIu2zIGwBKa46a37kROMDEQSG1BbmXvbaDcQ
eHRty22jV7hBHoy4GPnNWEGcum+cYr1MgxoKInsR7uTSClqwr51Cu9EnttICXd+F
LXxIL1tG95PCdHemv17A+ExCGllNMuDK79AG8ftd12s79M5Tyb0Eofwoxu1IBCTC
Iq0YZ3tU5EZpmqnyYknmnk7UlgiaczjFVZ0xd16ft1wRSM/00rxYyAxoDgo4g+y5
jjHSfP4zBQo+jijOpRINRhKGZy34rbzWIYQv+hRno9c9BKQbkirFTnVpTJ2k0xIr
bh8JvH+Y+pxll8BzzcKy64/FqJt6lGX0CApfP9vcO44eF2OFrDVj0DqFlvobf7nw
ReobyJA9KbHPlLwrjLv5KE26aBAWCEHNYvMD8k2UDeJ1gaHS03kmD2fa/joBjImz
iiHSi7mbbTWy1vTyKy47w3qV8QCQCJeZpArBhNM/3oPcQzPvv8PVv961/SdK3g8J
+jOW4aRbHbU5zgCBjr/laMBromQcaHcupTbK4yNLzzj5KfinRIZpOb/96rSh1X8P
HAI8Vgi8xUf2h+gdVpY0YySjPbuMO7fqdYnB7+j85LwlgGP78ceAaUCwjbcusg7j
FpBXNO9pyZUU1zG2DuMKYE4NCpP7KDZNbCPfnVMlP7SrFhnDNFtg8LLC0lAVOSzp
H2N0oR5zpuFZETqGwgyNAPJdbx3YmqsBEYPmTVVIQjcWyt4/lcAmAOjq3AoIIR0U
R84IrjS2t9R41sTUInpK4cFQ49RqaMijBmkX0vUTFUs5LTwXtK4JK1LXDjJp0/Sg
yhCfPWgj5mXbNgf5Lc2kBTJ9RWviPTwhVfUxmBKLH+7ArzsuIw7nO9IM1dWIRZvS
/35DaUeCJlULl6lX08+HYf1bmx9Wk0Tg/XigD8TicF4WuxTCaYkZSkvQlyu/1FCH
iuYdRzDQ3g8Y/NKW2+IStcGaIYAHlQBwr5hEVwh04EMdOsuw47WjOTl41DvrEA1a
Zuu6N7Cg7HoB5dyzw8pUmfzSwaVyyvgSkQ1tr2ufumBXy2KTN0IO0/h0F4+UzY9D
tQh44g+oDpaEhzUzyukScQb4h6CRGzsOtlHDuz7FzaFxG9B9oltk/IaCCQUQnwCX
T4RhScwswC3q0CL2yTY4FbvD7WLlzP1b19uA0V0GmRa9/5BMBYfmIynF36ejOhIc
pBZ59QwNeuwawAULo8BLqGqIMRhiu/u1f7zLfmVmdYLVNt7CfhepSWFJEoa0gbnc
U5Z4rDcO3iTFF3vsYwiGTmc6XplLw9yXz1tTBz5Fd3VQX5lwu3UbtptOgn/8hR/V
Y1jdeZSSLgcOO+XJ8NJqg3JXSrZ8ZDiPbvEu/lgitgcrc4csK5Yiy/Hn1XDjDD1l
f0BVdpD8ugjTnNQKbYutQCcM5oUwOZeJKo4D1a+4kP9E0/cjBdkDSHmMAStTUuBw
ig1QaqlTCNFgM1ruLy6BR8s8f24axkmkhlHnWDDCupdFDP211I6cTYgyMzgQhUmD
/2p0j9O3Ijs7iBE/38RA86KSwojcS1lxppM/sd+NzliTbqc4vNHj714coXfVIOWC
/fjNp8wJMREJqZaEy22MW7ds1zMTCInrQ8/6ui164KOOfKIjQH48C5uMreXYKtNb
HHsMdGD+8OnShtntqoK49xEAtYqKdbzNxh2Z5pTuVhUtAEdBZRXIKzoBZSPpsoHr
wJaqdSvYOMIFPQKCptCJMOc2Trtorprz6n1enTo825OtWdscLFBMEUoWP+MJo6sX
lvRAy236xyPyarM1IcS+Kss9ahSLdLsx1avRaET5dgC6l6aGtL6fq7fWzRmqKLsg
BJUx0SjJIpJmv/5TzOF++DXvIDAHIxDoWynUJrRVwkhR4Bj44dEQHziWIbkufQl+
QykkPvhrQmKPAcRjHz9JQYrFrxFMWJ0+CLTRvPhlATEvX6vQXLSW1sjAjhdcgeuU
oNUlXACl1ymNroa5aNzOMEO+1mTvpZCU7N62uVGe6ygAtf33WdAXZXHF/MqreK7x
fl+Sv4ESNDfx2nPJf9EuMxcuk34S0Y4yGmLT+UodPR0HFGHYk0KQGfGy3oc9ga1H
6NlmINn7+6ac5JXLAZPx/2fWuYyvpvIqzpANc46bKFxloTcpSs6G2wA102+3E+gD
Xjgtnsd9sH6UaK+7gWkpU+n3g7WIwKuNL/dvJa0/zpR9FJ2DAiZlxNvT8vbIWZv8
GCzZ9q+/93Ct9kkTSi86FOeGcWroCo9c4yxErsVwFkLaAEDWXYh8irUVQ7Z4BxQa
gv0a9Na2k7PTMLDAJRTbSuvxOya/4uOdFApeDraYdv7+St3OmimMPCb9wsEPAvo5
mypY1q0atbfXgj5Ng9onNesAYqZm8ZlCtehoxDtXSfuDiMjSh/4+CwdZQx3QUv3a
2jCrJnY1CYYuCdP7+FThG7IHjOG31uKnGIa5Ouw0vh1RCDX5TbW4ZxwltQffiqmL
4cOaPJ+ADD+BVO833ZHJjpnJrIZjLtQtXlFmze4PS1iBDZfqoKLlGE+m630Tcrk1
wPLObu+LLH4p2qxGkWAMkPe0ht3LKanhB+2clWpFAtesQb5w8ppUH4/L/45LTSLX
MMmqyZN+3pxOu/9cybRSOtbxHR5WmPvjK/5SdDHP13Em8lxMTbGrGgPg1rnQvmgF
Umo01zw0F8HqAavm84xK9lYMW8j7hQOd13EGJh3s2XLWCaiSzPbigdasy4EDACJg
PYIi5S9vavm99uY82DsWRMK50fpM6wvzByXRdqG0Np+swQAnWLZsy2gAuMJNWRHl
v1QQIYJGexdDswigwr1SuNetSWtNC3nNGrfNI8+FKCfcC+xbUCIZjnGWST97t+VK
/eyxC8qIrJpO0HF3MnWI31E7WAbGRcSO+fR5ISNWaT+EMya1IN/sQzhfnEQcHudW
hbkr+aF7LHvSrTlDsXcUrAVPCz7b6UqcSNi7RWZ2++UJQHZi8yxDXGizkc2HLX50
8JFlBgXOb+Hx1cCTDLnisASxZBi5EpnfY1UUXKbhJMYriBNO0jxcBMhbuqD1tmM+
JwVOCglqkyHwT6ln7P98KwQU6dHiB/7rZQsGLYjMcB2d6e9Pmso5sgcpxZCf3/wQ
mGtHUmjUm0GkXpNrD5Kg6m7BeDjqg2tDXhiOECzMp85rpI/YSE5R610k0APGhh3h
yB6MeCSAvOXKZ+h/6yubRfc7CodHLGDS8Uyu5f20hBxov+7r7/TOqpShGnJRwxl7
ZXf9LQ6682hjHrNLKX+YWX6X/YGQjEphKwTLW3do4Izs3dCaoTRlCmvLm2ltOSmi
7KegjQkG2lT2Kcy+v+haRsZHxUYYlPUp1USVplPlgeSQWfpKEImDYSBQnJ24zllB
+WHasseMBAdnqIVuH/2Qvcq47IV1h48uONE7jP+tG4DOfEAzEj8n0SF5IeAiu1+W
I5z3FGAix+HMNH4f6sOBudBEaP0ae4nXlmUXsTLu4spHaXHwOLyNoWiTAiEWj6p3
RaCLAj7Ed8THfrKaVNMVMzLWCetkUC1ujsTtFTPWPGMEActhzVN2MDq6sej3YiDB
cm/+jYaVwvF705VV+xl31+XAzmoTgrAI5xRRs/079lZqX25k1AjOxJXBtFCoQY9T
Gr0YxzqGDQwbG0RCWjZ7CSv+Ugn2hjPb6M635hvke8xHdZzGqxljks0e3k876z/e
gXCEpHP1wrNCqprOnG2jkeR0bmuH3w4+LS1MhaDyuj52oaHg7oE/Oz2LAlKNl6rE
Vgh3OEMCM0OKajCa+9xIQUi4al3jdRLqcauucYwi49PedV4kNzOTiBfJyKxpq3E6
EcYmmZmguejW4OM3FU0OBhyQBNDGUAZm2lNd1e0WwM9UfiLgNx+LwT0rNlwTHEDG
y6Q0u4XItbH//g2h5udfiWQKDDr00IB9XAKoOmbNIvvbzFOwdoNtiSHUI75ywCH2
OVfvNQUUXx5SJXE9Fs4B4eTThlSD1QNCGrE5EWif2pfakV94zaoyuKfObUHxeCuw
vAtR34WcHE7HLc1U54fX3jENf769GBBJNeFxT4aQIk1dHzxte+w8nhEI98WqXGGO
V6ThN7BdAc0jqx6+oDWDyvr/LpyV37FYCqNyhE860Ed+DCiM9P+wxHjV5wIgW/hF
Padhgsv4jou7zbg8jPY272Sif+uFIkSj6HeoMPgKmtlO0C04z/zyLzxdbyoWuy5K
h/Xd8UlpZZv7nf55+cSixdQqqg77VLqp7PuWKDqPehSHEe+SR0YHiFzashZ+JsSZ
ewfdNfegLGjRwf2fWbNLSd0EoBOu+14FTrn2VYUiBSMpIh1s3mxzGpZotqMOkqEZ
IhxAGMiMW+MF4votXWqZ0Dzs6oF9hZKGqwd7qifRvo/yiRVsNsGU5bamfGeFCKy4
w92AYqifP2AaawjQuyKApDaE007sIaInNQ/ywjLn387hWkIPyvV9n+EbQ1Jjsh1P
mPqVfv9Ib8EIMFrMf1NiWgLaIMOI0Xkb2YCthwW0QsthDApMSY1H4MOxVYoUnTc0
2R119qmaQqejXevu2V6q9viXkaVa2ScUyCF7Zg67HmXdE70gUWMWXdyp6+CXvQob
XOJTWWwcKy092phStAK7fYwIdlI2cy2mlKXYZwIcNMj5J7MRo85u/tQtpIvZqJgk
TAvxDxwaMU3Ef4t3tDlV0Ak+NCo0u7VDsxu2lGSdCdqMgBr9D0LzKj6pulV1y8es
U0x3VgwEPRcabKZF8nodVroeUyiJzAlTOHs4G44MdbtUszjr678E8urd7EhQ3PNM
RusdtMkfIFmH+/djipL7Ms6740o/F+3f4RGYFLQXYqZ9cyNmawcpYs2HKUVssSsg
mPgbcx9qJlWwvwZJbn6m9ieL6t7qWw0kh1kEG+ET4CmKjT+UcvwqBWkz0huVqHB9
vCV9JRpDgbpkAQyhTxuLRXEWjfTH3OzO1R3X2dK6yFYki7+ajcxzUIif16+HiitE
J7/kju5Uqy5LuuwdfgBivGO+vN9aUOwzowzErHDeqsvqzimVu4fSAjuox/eykCzc
+pA5+79j4rLv59btp51FDbxo6EHDHNJJGgmhGLyVsOJDVm914fZneK+qtHIcjoeT
7PsiyvZ+ohdFksscFXY9jmDk8QVIQQn5TXuMZYQVFc61900H3lGeZV/gorAfdPmS
0s4xzvUCK8fK4YJvDXTASPvzppeKbQKQt2s6n3JFGepKicB0SmNA/O9CREmbGlt9
70p6EBbOpZTNDdQGhlAuY7YXgi7ccLFDlw+wg5AqFGgAjzC43sbOpX3pRoGRXTlt
3/yjCX5ECwcUhvsuYw/yQxURrJB8YQ/idVzsr6VnFCLZVuY51fzLjHJ/+V7B4unz
Ug1FKjGY4ITIWRCPTRjV56xDjjE2wgao+Xmd3UTI08olf1npxKfqPohGyHsOrWRF
y4MpwzE/b4LdLeVSaUol96ggRhY8LDrBOYSfxcNt22bOqJTUgLazvfL4WmZo7jKy
SmU3BQg7//whjvQh/InOdOWWblyK1tJHX5/lIwjxPaUrXQ/GaGsjgnwy6jgwDF54
6BbHOvW5tn+HdJB7Pka/0Io63SVYaBttiW/0vV56h4Ck4usm0LwGaCID9il/LlcG
KEv9W6mU10a1nd729+b6AVgFMJw+ZakS+8U8ONgZPvW1B+Yqe/B7SWcCE9Pij0QX
uDL7uzPB3dEG3xYLSSR+aFTEjRl6fG4V5i0z+mKf4OwZWDi64kAm6BnXYT9905iG
7hG9jeJfmU/HOcx7TT+S6ipvKJX+Nzw6+6H/zirSrE7LoL1qDsnHNDKwIzFykbES
YB9qB+KEL8GmWPL1783hSaFHqW87RiAiwOZCUdw/8bW7Rk8JIRKWC8txmObPr/qa
ZOMZBY8gU5lvFLivMXma2Jy2UtSexwYOELQ6ky8wcUGeeexQXVI1kdWCuzxZozGe
P1SlGZ8TGUJ8uhNVfJMIB9vW+uMRqTzGVBLJ0pR/Sr8lclLZzW0E62fmmCQyqZ6Q
qfBQCnNrIhyDTqa70MLKsMxsCq4/dvP/VhywYo99czfTOXnSxFlBzTlFLRQv9Va3
nLM9FYPcmH4OCuIhtLYIRy/UwsnrvTZ1+dVl7wMYjka7j0cl82LrO0rdRcBeN4Gf
+W+qQ39LC94DECtzKrw0xKWx7ufwKBcr+w+QMEEmGIRbBd8kgSA5CkSyOAhb2yYu
napmtfcM2X1/hrS9b3oe/zRDRI7KW/yoiMP+TrQZmM1bmB/oxw2yDTuiRlH6jhp0
accTaiWpBe/MWseRHGGGxYXp7hnQmlemIO7nSJFcpD7EU4UDECcjS8JDDZa5Fo+r
cIbck5nFnTK8Jb2IEpnJkwzN5Q+EiLF9XHv++hzoDa/0HiQXCLTgAIZd7pwuXqDN
/4EY5XUyY79gW94QJKWGmPBca5fHMgCoe3JETmrcuAv+POYlKZNvuIIALVlaeW/E
Z7h7RE42Ze5e/8YFLsrx9aNJqHUNqIBCXbK9mCv4GjqVAKvXSf8HCbiTq66GUfJu
s5xqwVJWVNgnSFhKU6ULiFtPM6iSHoAMpudY5k7TdI1ppQrWyqPdRqSz486Yxhtr
ah+UQtB7eK0upKm95zb6UMQzI5aEm25cbZgyTDNtwF10npk3uayxHDqATj6HNNj8
EUQBP6AFPTnk7elr1Ip2N6YUt0ewi6IJPyUsrflxl+D0bEzGXoG8yPC4pNrSH2B5
WEaKKjPouHkG9I97CxViyrXLM3cJ81ycZjLwGICgs5T5uFMlAgVCH2JLPLdxT2l8
+hhH96nB7/ZQxa0PStDPpYmd4SFnlK/FlpVaWi9tLmA0NL5JD3v3fcqojcMDM0N0
BurTArAv92W36zjcCIT/8nuxuafM/ggxFq4MHfjQ03Iwt3vGF3iwi+wnA46pRlbV
RAbifdtere8T8jrN7iPI97kUfqiS5zECYD8SQpjP36ji8eLU7SWOmHnG0QKOgwRb
XJ0Kexj7L6CUqQKqlE+zXW3HGAzRlLBe2RPgmD6BqcgSJCunfYCSzvzqfTaNibT5
gqHpFxsXAy/8w+IrrQVvDzrl/ddyWie+uAXrg9q7rnOhH6JmQ1NVjE49xrgRmykC
PXaD35/foSoMLGRwNsopInBQdYFQuc1i5iTwOkx+G++WbzQxOJu0Lg4LFYKWxS+3
8+ah0fxPXDM9+6XHFeISImo2kSXXnG/upihD4EAceJeb3w4InMQhpojTHhZBOzSZ
ltCBhw9iI363vrF1wFIrRuCA0kWPkzued28t0E57sbZw59ogoEgwHimdiD2w/00w
hXCcTdqA+pwlR+IKc2IHV1JUcTwsb+ja3oYG3ouYQtQwbGXu50ZxSH5tVOI7q9+0
IbbWRn2ykITUAWQtJCWwW5UtpKNU8/fTIOWOOxf1rvOeuxJz06u4zDxIWgOLF7ut
BkZX3ooYRlLP8fqx446Ne6OixCsf4+RXbSDWyMbMA9+6KZyRQTAXmOkWQaFsJfOD
8vC4WCX3gmrO0hHl4q39cBr9ZqJ2wnb4CrX0L/ft4XtGCnr33ZgyPT7graDkTu2z
fqVo2NvcVkMFr4AlpxWrFIY5Svfys9dH+wK2qM7rS6gtETpkiecc4LFfMVGxP62l
EC6JIyvNUwdmcUtUCb+2TPBLR/kicyNJLYHop+hvqpzFtRXKJRVbfy50fIVMSNlh
gCOVSosd9hnGAilZj7uxuUJLTx++64+xqqhQ25v0UHC3P1rcEymLw6z/CfqJCe84
1Udx7QCHB9BNO3XDFnZ+jT6UzlqnTvt/Y/u05t6FwsJe7aYnpOrWnqRogJyDotna
sEOVgqnmEhc1BAaSE93/iyPlBDwj6pjwetL0hv82lApvKOkdN6DvOPpZB00RO8Pu
p6KrKVycTTYiqU3rFHNcm1XW2gMbC12ifBQ4JfA/utWIlYY4XRegkPTp8aEpavQz
7SNu7AOFmwrZ/iOlGSNrob8VCJ2HGpAe/avB/Y+1QpdPpC68RT0cPi0EDiarNAH7
DbjnADkcw2x14HSACoZ28ybJD4BkGGo6QX1/7OXneDuncv+YA6TQxDrW7Cl/hkce
wgtvFSb7ImvOS9MrR6chJhdGhEIR17B2HecltQGc2ykTsZ1YtQTKl2lOhbQuPr/q
UWbCFiazhoBMh6yZecFtCe3xJzp3VU347WK4dKWBMKkuTvk40PQmwTL7W+sIxH73
olMPp8R7/DuysFf4Gd5X7jmQ01+vauoigv3l71JHBEk8kIhtxPpKeiPyEEqwPCCu
9EmAiCPWsvvdJm3EtluiaeOHwLnK/Ani9KDjDex/5L87PtPLU83w4jL96eqEkuhr
7XKcobXn3bqB86G3kApZC1VGx4ZrKk96Xl+LJAD5R95njai2Yu8g+rKBtHruOCPY
2jtqKTkRU2A9fTALcVbxchNVp8BCbbOj/8M0DgRxSh8VU40eNSZsm/CfdWfcLmng
tSdpUEK2ExIyxOaNoJwRgd/Y5dPFW1DmnCaL9xMtTNWiJWB+pdoDnDnpICb2GbF3
bM2t1bdOYOVGN+sevZqGeaZRC/WI1mRf9nplltIKezVX8ofaFP+2010IrZD2GHUm
uTl+8DV1tYnxgmbjvW9aOXJoHieOteNe6BIQEb0WWxxrJnxvtS54Gq5zQqpgew2M
bkH89LWvz6n7jzFDLYLzR8Dugx0DcHJXIozCP4ryZRIG9TIb6SXF5Zc7AQ+ZOmbE
M/wfctDjkm+UCN8U5C80X/Fs9s6tyfJNQotwZeGS68OJQ5ztSit6Acv1jU4CAlAB
WNRoknQ2X0c/S6my/w42DLpGu9o2y4p4WILmV1B0X9ulsfIcX4HbAaNrPQsp7yP5
Yny2iCUDMVSETUxdUdmLbGzHfQpsYxz86YulRsdJtCg3+ZZ0c8We7NGBLCFk/86E
7ETZH//60YyXVDuXMIqfDfRRQwfQqWdsGQRxFAz6Po9SOwzEA6FUyekp053E35TB
oRvspTSN95RWfCbT7vkQzgX2LGkJqU6W1d7ZX49DqUh8MA43QAm24Y9unSib5MNW
En0NCaI87mF+M3PZQYcV7kIBIenP6IJtoG7paAKzmxEnpFCkjCi6nhsTdJJ0SoOD
ji2hqOEThpw8cfjdT7dnoglQa0b6w7zJgmdQqIk323rFl3PR5D5eZmgItpjQz+sH
I9Uv4GIXafl+EHKP4v1Cm871Oo/lLbPN6Iqq8PLGxtzNlOXFYEX8BKaGn7lTApaf
aOF8rF2vNLUlaPgTxzrjB0Mi5VMIbVCVz063o1cdZlnwHyyBGr+4FtAnZA0NGPkR
SXdHO5ezlMWMlXyWBczgdnUArltFqlIyCSNeYPtBMysWlckmlFNBJNKvjA/5Hbm4
NDex5aaQc/Qg0LDbRCNKD/zQXMlFT9UzVP14tcYdodNel7IUgMNHApuKrqso/1t7
vckdaxsjgwYCY/oTJxQTrihlsn8UlWasitgn3ECJiFCKYEotqzyesWmbMxbunjbN
KQkT87dYVOWvhYXuy8vmqq+G+yIoj3yYt7EeMRPOUSp9EV5X+oBgyetrYZxAZO5q
ztjcPPw7j28M6vO2M7/ho8irv02BaQpd7yPusa2YpREMVSE0oKB1OmePCceFuJJ6
6faYEQTkivFP4oxY2SUb1ssKlcTISOWLMfmLtBAyTPaRdEqiRNXgFtmZ31WedXCh
n5zi8AcQpLkMaoRiikGFvNEzz2DVtoCz8VfVNZmapI4iNe3LUni6R5nQINqc333I
tiRW6eGto46RAgShVTD3Y8rpPrVe46Rf58izEsiWIaGVM7njgYykmFz8foTGa1dX
fJWu8XLYIuwzAeuuSGKJ57WNmtZg/Bld61CNc9bTrt2WyqG3Ov23xZvbcul1k5A7
T6GutdLzV764lJ347wddIeuv+dETkt5ZVIrJQjTYV8gy+LlbkrNyfzqLDqCFTHIR
S3DBpfHPru5C2thaHcJn3Vi4fxfj81BH6yOgANtvxMhNWxok8LfLI99JXrCNJ/84
kvUO5L8ByeTt9vRhDymTRhNfNANHXp7YdunyHJbXEsjtjVH45+RDxRBmDLzcCkzS
z5lsqR1lDTB5s664CUhP89/5bdDdC0cAUM+C59o/FH4aVRao4Oqfh1rurexQZFXW
YNQ5u+G0JCYl/gja36KZ3T1KMAJQnCTzsZNk1XCmcaUAikCC4JIEmzF/F9lqPR+T
0kPxEWD3wpsjSDVtXII1x9XhDsuaJ+mkqi5bH0PZbS+ABr+HPK8W08vf5TF91tHL
89rVJTylXpow4f4gjI7Fq1Wf4ajZN7aGn4qBr4nJQNpM60xrca/UzocanUqID35I
LoWB9Qk/5T/y+UQOhF77vFOc9IP1lXW+lpGD/+TCWYbZ+ZcMsypjA1cnrZfXv4r+
uW1SaJ42Ay+9nDsjlqEK4+lzMH2HATOxaE09g2Br6BQF1WHk3Gi9QS4vGlpciRe6
NjtGfCX4PnqlDLnPejKcT/PZ1rqz9e8Z3hDuwVebLIPOIO/+YOJ0yDrOTKKhCxNe
JSkSIhDguuOiWmpEDwxvyi9uWO5PL6wIUQ8FZrJvoZURrmN28ZBCanuRtydAeMyu
qkrDhjmK3tQD4VLPPrcgpUhRbS3Sb44/ApXJPFpg7e5OL5nD/YqDjWVFttfqrXsh
tpj2iJLajY88/iApekAvqtq+Qktrd/99HdO1Bg160IA2Bjet6UMP+dRr6UPrErh3
/RTCxGulyjp3LYMBfhgmnOnM8cQbo7J57X9kmEtxTzIpR4QXTm+KBfvwyFKYY/xu
tn4DLNzgi8nhh7yIvBD46V8DpXFMTPB6I6C05nouwXjPjGLcmZszYLPwgnzOomFf
cqOHZB4EwyPoax2eJqxnKjOw6dpL7alIpeJE3fXaugiGU/RVvL97e7vymebIEqd+
0UJY4RV0COeqJo86BknfIiUeHhgEPgYQ2qW/xTcy+E6jswb7a3Vt67RPECMav0G4
yzo0GUG1VyF0KSczUIsyd3bFonW428z3qqgDzkmC5hgAJkN8OKo0VSja49GnPlbo
rxa2dr2UKp8aPMceySAz7BKpRDnt/ftBBiYS6MwZq2o0NF5Uk47OgzarPKC0h8WP
6tyEA9irmKJJxrsoQZdNlbsk3dl/ve3FY+Mfexpud5IpdyG6vqqeLTAlR0bIXWTl
LrZktrp3Od0MQkMYqwJMPYg7+MoYtDICkj4fQ9Zpm7zm43cV4DL56AQIbT2g7CYp
sXpfJDexXKEHLhddtesxXJw1Pe5XjY6hnRRWpZHMyOdMYkYW/C+LcOg8rKU4kasp
lfP5448j8PTsD1yj8kXiYD4Bwq9dLJEFqfoORtHtAsxQ9CYmjlEKUdvPCvn6B3TL
hckEPV7Yop/dQkbuF8doadw7xMj8AUGgFCZ1T9sS0G+lQtFx9La49q3FsK0Jqd9d
cxQ6NNAqo2xPBR7Vq9w3FTGMf9JTYWQvBhAItMJ7tnulCeKMfZY4b0R5yq6euUkl
zGzV8I0wVE1RZ6vFD4XTTZ5EkKC/AdMLtZNXEnS3XlLhikBEPBjbUhkdNKNFyWoU
brz1Rna6RuqHDRh9LANkP9u1O9MPQQiItSP3TGF35EqhBcRNThmHRNjohuuMDaGc
MVEstSIUzTxNH7nOyCmParDOGZp5YGn2K7niUdlXnUtYlCU2RBkL0otBc+Qo4LHX
8yxcYhQCCz6cxUAAiPvUpvwo2WV11LMp9ULpguvoqXhj+xk5lTbnBntmbrxUCKdg
HAYvCMnJUxjFgMGLYi7kELwBG1r+x0VvRjy8dpGzOb1a57dX0pC3IXsEBtvSnehX
pV1BGDhwaEWyxXg/4F7JCiZxLLojsi6w8y3wEf/TRAHd8PElSCOU+MEn01eDUBm7
90PWPSLo8dzQKyctxDLhreEtjImfUvqbRUWR21swkOAsPOlh8UHzNePljQh0c99W
sfv4sTwLna16RcYZQAAUwjQesYtfgUMRkUpKk6dLAEDNSEUBxPzskq0IRF+0Ycf1
4/UXo9BNYqdhQdIACZ6uc5YFkGml/Z1STGze8OT33yk6C0j7l9MwahJzmWDql5UI
ry7BXG0WgT6SCYJD/HLKm0f//Pa2A61ISlu+KIkXvf4FBKTdGeNh/JfbYeCzwfla
mzZ/H4ZIuGHyqMsaeGhhWiOfBDddlV5O7nV/Fa622FcKcqgd1HwEMgEfc18nGDqd
J7zPsGaxRejSnIqo3Vv9QgJiKQghXypavUC7NOKakdIL0Lndq3cpZ7aG0pE/OrKj
RgMaOQ9loJOK0Z0+lnDdYAGVaKy5vomBkVjsVT/nBr0CNHvINKosQwMo1dyM6xFb
4jeNlNC3U1jf9+kskQj9zmWQ2ZFVUNWXKWP9lu1iePvkbKmnZ2ziAmFR+WIbixRd
YB1fch6fsy9HSAuV80LueNRhPLpl0/Me9/Tuhu2cEmnZdJ5/3T3yQjUGK8FgXraF
dw8w17cFXErJifqwuTLPf//Rl9Zns3oGlTdACLvFkym7CMuar/4z8TVn4Ks712Mj
VY0JhbgYunKt3B6TSlNfBxUUYY4NM+PqJHJr6dE/PYEh3wSPFIbdaLxmAdWplNqb
ZcKORhGhrPggGb0Y6U+Z6Sf11GGmyj8uzbNqxOcR13F8TDvVALcpzA2UYXESPyEy
UjowyueWB5a3+nT3uY3UizeGSsS0qiIr4WIDZ1XCZUDLY5GPE2xQ+Mk9wkH6q7k4
wY7/QR8/NgvAMPzRz5xvmLU/USnMwsjciFsmIRTbT2KJky4oSnTQqHx2vl7frGFi
yBX+mHpUM0uDJKnOernw9V7F3vjMoBWd4m6TVv/eMCGcz8D9vgLMQv6tWyhEUwjj
bx90JCvnYgfHfoTWHziV7MNRIviZGXRUGRCzwWmiBHcRey6qmoHGAn2akC4uFmCn
lB/xls1aW2J3mRXApqN8YUaugu34XqQ9C3N3GKY4nJLLEQhh+Ptezk9A2dbjbryu
IfgNM3wCCJX3YvNwKxc0guprnvjhG3YfklyxhzMJzlQqXC0OzUQ3UQqsOPi2AjNZ
LppkbRJe8TRLFr7JV99oxCkGRnKgB9uDbjam5vVcWVvNC2RWeRFWzBVJEnqVKOy5
PSE+c7VgKkCvWW4g96eMhFZ8Rtq4JbDvngtATUqxPCM1kLJQNdwTOwFpqjIVc1+u
jZBnjxlk1BeiwF7gnPYPBdpUl2SOKrbzfzQID34UP4WJhd24bD4PuQ60Ew1yjVAA
mFySI7ynajGr2DLb78BobM8X/SGJAjCvL8G+gqx1tTwywE4kY554uOikIznQnRNC
o3IzlYp/7py6530emjQ5u6LggxyjO8B9a8og7jG7AQUJh1rmfHkLWnPWji62jMRL
5/8LTh4iP0efzVdZhyMCx+IfoJAhe9+6b2/jck/rWIFNg8zyWc0cDf7aXapnToY9
z5Zh2K6PJ5Zekqt4L7Tj92q+zBDlfFK+EfHTYYs401SzI1vKJlaugCLnwJqy3gcf
zOuqnSZGlXJxwWVVWizWezPczLs0GQ6uG4ZJpKSg1Cpxm0SXadadNkKjnvd9ry4a
oKiasxUim4xvvesncoic4fuyFKo6s9OplpqopJXgvFA624p9MPl6s5oz4ANBN5I6
kuezGSMnRktozqoZeSL3T12v0Anf9maeCjA2hSkecQsuJaqo1cS881Voclbr6aKx
6bjnsOUIUcI/QTmcLGIZNUyeo6nEa++PPdJkIEzkdITkDEEOij9kNBPtb9D84laa
i1Bar2evVsK9npaRWVOKwlnpdhPhRW4cPCgXpkptlE5iphOxLKE0RW2p3PCJin12
EXyPV9dKqA9hqNoJPLYDHjdKNRh9XTb+HvLeyA+dsLcMf9zOpftEHeB+lrV/7+VP
OZk0wDWCTy/C0wf7MxHf+tdbYWNS0Oqy/yhG0wc2gIw7yPdADbUJO0gQhFviO3ic
hFFcj2FHOU8SH2r2jNWLyaCpougzP9nVath8ZleNRMGDQ1e25yp2GXACHajgDzSO
79FMzZ3rCOmZOCGE9VswYF8YmMfPxyHAtsRxQHLgvJPluIZqNpjonB+IMoV2xMt1
FAQqPOQCjePabXrU1RlyDayANcF40RpERf9delMSDd6HKtQ9dvONF0bML/jG0QVf
GNV6/Ih0DrWeuZl81rU5B2tvb79sesyukoouGBvtY298RE0Zw52W1mx9dzhaQLCx
9SaEZomDSzmeuwvx+8kqsh6zKMsEx9UdbgxCeFPZ4ph2kV8roR3dGQI8jgDfleuQ
RLaZ3BSxgKumDr+tILiDWlUf4+jNm7NxNhC1l2rSixjLu5LzZWOrQCEBPWnC3Pko
0bTwNHqksJYzNCNke1kY5vH1EgSRY2RIKJPFsvQL06AXF4YSLOMfuB6P6pCAna5y
lnkF6qB5lV8Uw3kpsQL0G9++2DxaJwAnthi0ouYa/cxDKH8TF6vVt0n1qI9+MBoZ
m8e/f63rYYV5v1rZEfvTch5XO9Ix2+VPERulVAD6swgG9JTEIBtQZ6FdaZ7p/zUf
Qgtampx/xKLTBFQJAijasA4OaFM0qk9/331KoXizxoR5xzv8Zo8WwrXGzsFgV8vV
dsRuUUaUchqeAd+igLN4GZjCLGXf8v9eTY/ByZqnLlnmTWSAKByV86M/7jC+lwam
M/ITbKqdQxrVGCVW9E5i6qaDXcvTv7r5bIT19t0r5CvLRf4DxNkm9WGEwRsfSapM
ddbk85IxDwiIL+r9dn1vblAu6K7vVR61A3EF+6LSjQW4d4n6/o90s9DQgDK5GVUw
qTAFrP0YFIN7jNLxhQ7WhQf9jbPGjV7kxzTthRoFKbvXMCRsshG5M1V7gavyyKnL
bpPmeEu+copn89xvpURtKtE5zot6Xx+OBsEtd7Mn0ZOrVoLBeeVKVwcuOKdV15IP
hK6mMz19F714jeonqN5dXg==
`pragma protect end_protected
