// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:39 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YSnlpkez3UcbMX9ePDWj2vMmo91gm08IwFdYyiI0A+tXJR0cxcDZXb3XHLJHeTey
Dds/VDqbRO9VMlOSVWI5WfzqXKPN6NtXa49jDFBOLSor8s4SqaYevggWH8ljdNYB
K1aEaImx5SqaoygiwDiuhkBtNJa9Kzvh4zdGHeWkI1c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4864)
4dNr7XeLJgzu2b7lqJ7dlKSKAkYE6lEhQ+cqyJlZpxo4kqE7O6yP3+2JKsfUeHrm
/L+ZWjoMYlYqxDKZ9MiEngxh7ybzGqzKatwferMYqYjcw78j4XZg01MAObnC6HlY
Rtl2CLDJltFmeUeLOGUJ1h1FOaTbWl5XH24yv+VtzH5hq6D3YZrhhqb7ySi0Mi4G
5WVcUWinzPhRSN27IJZSPWAW8CfGm0IBBK8vq1rGfI8b+l5X1iVtsi9tcCQpKr+u
rpZZGH+mZQ6HtSPdVdkOm9DzjMP0MZCct0GMcSvSnXDjrOTiFGyHC36Y2Vb67yo6
2eNY0qFwPtBs0ftLlCGfD+fTuLJ/RSkRLxLuq2yoQdBjKWjajAsH9mo1J1nKbgj9
prEGrz44tGTjdOmAn0IRItlp9s4aaOUKp+pQAuDDbUcQJbDMkhowgYzpUaNWX5Sw
NL/MmN4f8EYnPd/eQo6sKWbGASm1UYALdYxd+5H7gi+p0czeNVv6ZN43f1uB3/Bu
RdbdVDCiiBgIm2KC/nl/GNy9d+UM2DLn0U5SMA4LUjz5BUPEUoLfbFjdp4azY27b
h6ySYkO9f3SVsJ7E3q1DIilR5tV1wZpSm0yuZ6VLwtMF3N/F1XcTlsGcKinMKfUn
p1fqypwi6qxjBHH/nc395GGKSTMivD5NYRpRQtFRHniJQVYnCor8j3kCKk1sd5BG
TWRUibguLyoyxVO8FxapjtLJGAKnSa2T34VYCuXTfx381wcoqSN4Crg/5n8yLXrT
wfTCz8LldM6qKgHNVB2j2ogAODx85FQIzWrQqAjjfsxJOOVbLlxDEMHsD+rFcnY3
ZI40zPoBJo30SwQA3qBJzUpE8jPP8rtzCyiCmPSkTzsxXLFfLW7eDxKxqMb7kW7l
ImCkxGIow7bKWXOtSNtva65JaMy6b8sZToyYDtFb+AdNa81ddlXucanugBSxw36D
fBX/nGxgnhVwomhfrhVNWjzSq8DYO1uitapjf9wZGkeG0DsN9CBSLzLXwaM/Tmu0
CbQkXxcO7lOoYiVYCv+Szt9wVO3S936B0HhvJsX0CXM7++RpSpEbxt9onytIrlte
cL1dnBCiMy+EfR1wQIaOb7lAvb0G7btoZl8C/QplpmEbA9MeT0g0aC2obXvpmwK+
5mfX+iZkzzdV1auGOVQAh0i3L2+FWre0mWcdzWT0h3id3/32kJWeSfs8kxXEC0xR
0Ei+VRAwUz+cb3xcd+Jq91XsGLAdHygU/paZXMiDioO70QKQPCXPokKIsIzl5F8o
PyOhPOFSIA6ByBS07+8Idi6cHKb+/VamIbExXSio3wHwL94/keT/+9NAKXod6ivr
CPDtW3EwxLO63U6/Xqa3TOX4d4QyI8K8iVPcAS6FvGpFuoAbNVYZ+0DFdH735zFM
f7I0hQAHh0z9/gED4NPZalQAVkH33E/LqQJHAjv+BRDzjDah5Fj2MuK3JvE4X43e
75vRaOK3Mr61zHpmbXd4ThZO+r0Q3tnGTJin7wHlzxollE4EmcFNG8ZhnOFMTYnJ
IJ74o0knNQoqbA3TrVuiur0AIt2bO38euwQK8fD8FgIYVuNhQYXGQp5z8mBrkCAW
MDY4jF+eFImYPp0l7i777zQApZ5mcyt3efEjCf1DpADcBdFJgXY9T84pA326JyWd
VRwT6euj35wMlCeqv8yStBCRaV4rTDT7I+qAy1RQERf2tPLXpk/HFtm7nm98/Ws6
S9nn8ZqRR6X3OzyAvbmVO3s+DVVKzngNvCVE3ULg4q7+jj02KnhVC9MJwiQe+Vae
vANMQ08mUux4Js0dHr6CXRw4BdvY93TcpV3JhBmDqthU2oZv/bFuawbnwPTLLf2/
78Ot8Mi1YFPLN967MRV5tLX0PPe+yVVpcPcNB9SL01urLL4xB9XHTDqCG3D9JQjI
ugYwlPSck4129TSetZ62BIhFhZZwutblvq3oS2Va7WOLheS2j9s9vaMwr4E8/x35
pFBpgs05+9uan3eutqi28OekLCOKEP95Urfg9evviXWrkbZtY4WD0uDiWZHnCZcn
xjwSHYRz/z3RQ2flHTfc8xRgPSyqT+YQ3cZTGszFWJlid6UZjI+O2sRP3dpxMAE0
UvPxrjdQESso1fWTnKmg0w4J0nJ9hLKF1gm3La40T74Y9sJsrbbxIV+vjYawRDzL
VfDRKoWZbT2fE2HssqjXqQm5EM82eAYdxIcEjUed9OGXr1YV7u260id4tNJhIaV1
FeRwyMU93jRhVWPyFqiWlLNXBVqCIa9H06qiotuw6CelU4yAswdTgjxM+KQ3mSqb
EzwSVz95P1VC1nqzyPwpYKtEzkUjv1YWOo1no6T7NLQ18Za/RJ1gYqCoLD+1biCn
JDEaeVgqVVsJlGyIq2BEmy+Caml9WUIldZTWr1NAp1553crYtpGyQMPI3TYGWcfn
I42vnkSvOeBMBhGDNyieqAPmthur54WJ4wUmWjow7UDYs/SiSxCboxqGjEeaOt9W
x4U1BlN9b1nvgLF051qmlz2zW4OwNV60DSal3Wth28o9PUsKzHVq3EznT2LnXVfo
Fw8PBg1E0C1cKVqD/sBcX8gcwKjt75wLcgNxpdlkdM/0q7lKTFDEDV9AK1iVq9I4
e7M3teeLQ53MYthUwibKVThNrJjy1sVnm8qz7H673MJwsFrgLpiss2kxzt4/70om
rvIM3PMW72TWKdbHOBdyTcAWBv12+m1jXuYh8LcaP2jPmJlfCyJ+fAapTQKVwcvk
F2HjBQ46D3qSlUtUJtL3pDiQ1hEoQCgCKhSxLjJvIVMVBDuNkd2LaPT2b0MFAOQ+
ZaQTS8H/ZNVdY1VCCr+UvU9jVJjFkAXR5/L5fvlC+F/NkAnJuZHiCCNNS14NQYLQ
cnhAD0te7TS25RBzPesWYlTGdaUHD0Y951xih8JSEaa7yvx9ldq50wzTkiZmDg9z
XmiF/5nHfxRmhDeVrI54GxvvKr7IzXdzreZIP9BXvy8NT0bXSYliz5QSs/yKLNXm
8bKfbKZlDIy3C5hxS5TWM8Qd7OWwpNs3fq/jwxzg7o2cDtcetzIkv+4qDRCgGY9G
TUqXVTJqOj0uUzzLfAPXhhhlsdy54vi9gnWPqTuXUiPe5zY3MfJpN+68BknPbpkg
5i14ySqqHl4JRCEpMFUMWLDVODktSJykEs0+u/yYVCUDdoIZtnSZccYvaDZh+lib
ibi3ne/X30Uc26f7NkVB8NioVZKVe+lJfgVWUTRZYtba0Z0E1L/UGJkpaMrGeZXd
ypmfQb3uVMxexTfVKWupLCOGu9cSkC0lNE+IOxMebrGSSbD9tzYquGJa/XOlr6Ot
T8n5o+M54G503mCtU+0suf78IlNLqRyT+YpqiyimjRcm537OogZB0+2iIWylHlvB
pzRxZNSu2PYwDpgApr6UgcXxfZUUYQMARYdaKUce+/ZD2A0oTnJClJtsxU/zNtXt
8h+6oc7BZNX5l6BlCz02JlNTXgY3VK9agbOAi2Ufa02ioBjrXECvZXbhrUGqGYbh
1LrPwLscONNjzMT193HXcCH3NK716v2IgNmhpWGNeSyUC70khZt9aVXVd6wsYlVZ
sXOFkchPkTGajeOl+c3Ubs4CWLAE3zU4VLwyh1BHTExN7Vvz86f6zsOJOuxLEDvT
xtr6McaGJ6hv/VsF+4fquRcfIkdx2ch4tpUkmB66cdR+5yz2gEANoas6d6yMFH4X
mymsK6+12bKHpjgDKH3ZKGIE+O2MrBaZ6n+Sz6Upsh1XZzOLjuKbwfqkIz4n+X4L
6gtvrtDs1q7dQuLDgG36+ocN+RIzgvhBThPslnsKKOxViI9p86REH0gW2RTVhKL3
2LF47RaWTc8TAJLQZPVquIMlzHTaoPbEn0DO2v1iggM4Gq41L+pP4ed5ewblvjIN
5X1WGdAIIpct89WpjAwqrGo+/RD/vvoaIHZkcTd08D1Ya4Cttz9yKBBA0cV5HSun
DUP8euEsY/n37e/TCwoqA7E+1j1QNa6F4BoWoaLGwraua0eiTT8p6Nw0CFc0XG/Y
O2bYp7d7NziuPBRaYIYwpdVFHr4suzGRODFQURDh3TvQgGMdC3xjB8YQ2aZpSg3K
kd7gSa2N9Tf4DSex4v7whhtuAcEhCiWMOLJ7/7W9OBu7VHFT2ABF+srtsvkrUZAG
cKrJtqxO2wALCumU0tMM7/qCa/K7mE8vEGH230JHWXRYisNGcctQp6RksctKDDZj
i44HXiHM1vPFuPtE6FXzCCphGcjig7N8OMnaCwL7WauDCewQjaoX8hBcbOmvUIgQ
a3CLI3AzbtODkbdtV8I74zJ3TvbOQKCThmUPumaxgFo2vhZmqnKFFnHatEhKjKi+
v8q7TuLWB5P0jK9VjG2YgoAKbG866VQBWfFffddOukC/8JCzuS2vttxTpfXjKDRH
vAmDIR+pndnlkkpCl6p7wBLAVYu0oWkWownQufctngHH3s4U3O3R5CTwmX4wvzWw
0//HdH4TsTHsTwUMSI0TfTIO1idddslbaKqIlRYFLkumMUzO8UI2z7BrFzJeKnvb
+1DA4MZTdmto36kroLiOgog+N6zP1ZjtYqREr0nWSA5zqfQB1I2pfNMNLPunKp5y
evv0ofQB4/a2jB8Mg8nPMjFbmT7ZKibedQNSe0HOH5mLnszBvZVr/7RyrW5vUjmj
Affr4wkiqilWE6CGCj4a2yyr2nAUGV+O4ul49PFvuI1cgQHiHJw2+LrcEtqDKhYQ
az1wAgnhY/4N0n4wLcqEU7rLQNxk7XUkK0q1O3AYtMSC8nxtBfnuM9tW+LHSKYEo
lU/ohuBMC8k0zK+1T4wNwFGS/Hz+sT/TbNKYPz+jI/iSiAFRWe5BzOuxFd5MAZgU
gowH5A3sVMXNdhp7G22nsgNFCv8tloQceC+tLMuq+aOhyUH11MmducOp7HKefHbA
OqxGCDwlphCYhnqjkJebTKEFBsfMHK/Acnoqpk/TsNXj5K09BqX7faqpRADQr1M9
ZXxuv8btlLVgzaHp47Eev+YyFjgcu1kmrZTusxwSfLUgElpsmra5EBhGSUuA52Xk
dGrrl5Ii/Whz215w9YNVPchV0Dx2eKSkE7fvYugPc7NynL1gK+rfVv3XwI3LunLd
fEnjGZdkipIqBOoZmSzDvO00x6C/DygFuSkqIAFfIMwWmxtmwofjp5WgJaBo2Tut
0/QyK03BBSzxLxsNT2Tju56alh1OYIAmmkTmu0sx49VRCsqWhlKqAPUC7AxsFs6/
oM3BEwTC7bDmaxTAydBXq/A1nkTpTtIWsOP4iOlUXdVMfxzvZ2ezX3+Moy3+75Rk
ONX+XbY9BaHkP2q03CXUbudD8MK5GneJDV06eiq5q6pey7BranDErlCIb6+PLcoi
QpeVI6KYj+ZOcR/tZcoXwCcinSlOrv2sJRRlqijIJnWWMBSqv56Ml3O6htDxCEai
dAknfp81u5xS6mWsuMuIGpYo3jBb/eEK1lGZWbrbDXMx6JivbIZoF3lWdfaGI39n
VKwz5ma6AiC2ZZSJtDHpF1f16GQyvNTubKMdM1X1AYec0f8dA/GG2yulZ+r8aKDB
H6tCIjhEI/EBuAsnV4r97xZ+MpCwayXtyXSv9J56/r6gnPj472oq88FaK8eCc1NV
3ZaGeupSJ3dgurnM6LktZpxQc5jG7HWf4iUbzXKr42G8xNaz4w2R7HdWoYylqcw+
EYlLCGga/G/KE1SqRKAeYKAR+4m5gzAG3/mDdsKCy95BzAnZajzPPMpPNFfvJjtx
ReARVVHXMpdujCD7X7LNLcOxpvow3wTcMCoVx7CJjoYPVR8mt9UujyWNjW+1Chdv
f7Oxe+s0yOjs2nRtbwylST29pi1uYKbDdB67FyzmgFxHYZXvRh6XE5KFivjULFZT
39tOQNEZMf53Ivu3dmiDJHdMLwSIECJDxEuBFc8Lufw5Xa6HSCwrZg8vW2lEoT19
vmG/BU36uOJRogaHJE0+YiY12aJgv/zH9EloKk/4pxItgsKWlgTfQCf3BdZjahm1
iQn8e2qJnBJ20tNODEarnmVsRyRlDJ4Dk0RpEttCQVh573MW07Orr4Fel4Zjjmrn
gIwxFkColq1eltAlnUGDdUyGlTaLvDjSMCmAv0uEm9c1fKoLLQvYu1YqZwWHuj32
6Zgc8dxnWUfKUAF0E8l08lYDLKl6N/B7ty+npYM4dwoTRlUi1PejiBPWNWhLEWiI
ZE/UyU3BX7sM2RTd7UPS3YJS7GQIle+NVRwIG4QspSjuA2914T1amEai9oL59DsW
9cgB/R2gtMi1isGx9d1TKx07ncGuAeeHg6mzw3zCjnKZsJ7G9kUrsZIdud0abSx3
6ms5U3FzAoTeL0sq2mlnJUFXGIHWh5carbu0QDW6qvjVFfv1Wki/EolwTmZBR2Oj
oaaPSa5kOFwAxYW8EsjXDi/q5yysLA6bh7osNH7EuEDAnjtl00Scw98XV2zZ2JCU
6MqX4E1hgTZ3shx2xakiCw==
`pragma protect end_protected
