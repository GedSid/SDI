// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:35 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cjtlXfp81H2XnIPwKae69AiwuLJsiGd8/T4bq+7rxyZwuTae+tkjI8jYeQ85CoKo
E1m2nes325GcCc6FnxkdwMHl45Vkiu/Tan97wBcJSe3ZcNQCp/Zsqa8Ua23vrRJ3
LSdYI28aWvVL3/03OBHx2rUop229hgqb8GDvPlDx9fg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 71104)
UFASACECFHsokXNwhaS74jD7Ewa1zr9f4cGev3v0p6JmT/MM5VHyMG2wIvKUNLu7
tlU5zrXreFge/JpZ5pBzOSQNP1g4UKgeZQjg/MYAwXq9aWqHLMRRDxCNC0/PBWjc
7zMBHwVXaq+bwLCuiu+iZs6mQnXXHixGHYhU+uRKdFMQLSHVHydBof8KPBso61L/
HiqB8ydGd+XT6/fCB8Zxtr6mHFYhB+eCUhlmpvl02uJCmbp4FM8QgdJ3tmKxNyx5
qVcI/e5WBhaQkDz8f9K6Bw0Hbn7JVt3yl4K1D6UzVvRbAWx8SM92XzQlFBFqmE+A
2Hks6tU+GsqnCbEF4u45QmeivYbsdpCB3DOgs3txdYIePuKINJtQwcEgepK+g02H
t37+AsCvF52w0lffToi1BE1kWdKohYLuEubIju4sx/vORIS1wxHakJZRx3Cx87ff
XJRcBykJOw8EE1KqMaL2WLYwZTvCC9ATOmm1YmmwchGkL14hnz55C56TxwFFnxou
CzPq7N2u9PLAqlVLQ+8b2QR27RWMxROw+ROYEddpzl8xOcfLhv+Rn+KCfphSpvon
HhduCtI7p5QLux4jkNXFPEf0jiSEKcjb+HZ+tFZgRkmP/KVNOhZPUSIjQCFhwFfR
QZ+mutfpmkm6Jx0F/Dne1DOTaa970U6h0viutaYt/LnmFp7r5BmCnGphJMW08FhX
1Js3dFFGnSDw+HwNXcA19YKoPo+Dd28/Xs4zag6tyECJgEqGrw8aXZC5wGMzThvi
JuF8vBUg+UIlKFT/fteCLMS5hK3Kla+bCg5mv9JEdundKQPSqSGB/sH4paK1xo6o
fouO8KnvVtSlc36l5o6aoXFAmvWkKMV0Shbx7XUnDthciVSWtOSBeQmrLEkZgk2p
vMunxeb1uUeLlyJ0Dk/cbkbuMHA1OmtW0Fie2rmFgJszfRH8oOkCcAwpiTWyqEES
Kw7ZEg358sdaCGGWzjAr1WKUckhlwDBkrwKDF9JixV2pSTkg4S4oWSSc1cdbQ+tB
aQwh19/KnuYItZKU8zWvRnrf537lXl3lF19OB559T0yYqXYPrFe4XTE7CX/auCPO
cLq8RiCdb/Ra2UtO5bwcLZ+m74VPj3zFbkuslaaPCECpupw+T2POe1OTJJN2vvMt
6KZYvAAoxd+5XnsWDJywaOLB8iMYU8qQdhvqzsZm5EdHfyzFMLmTSVgFvOceA9X/
WfiZFyEAse4bwt4RFNPDtiulZh45rGGKbkl4yflcn6/nPjiBToOWyS9c/sXi4KIY
/ey3aX9763rAM5mXFbWSDjHt2/0MVgjpEFqFmJ/3MHX61DoDOrRH6xgQu1N9vFDi
xhBxgWhAtqv95SWZ8w3C0OCQLiOuEWJVKslXX1inOvSFvHGUjXuaWpsrQhehycG8
ttkslGVTG5n+JpR/FoDzbSV6/0sxrNyatA4/BA4JlBpU3nVRbf3kK8yVQ+83gIz4
xrwJc2nxsXMFLdWwAgQHc6BAWpx50GrM/WHIpvWWbFCuN5h3wMXre//7P09EmgfH
r67y54fV4av3A+4Dv4UyZsK3iqyciPe5f/0xuBpkLKvRxf+XolMZq89qPsf/bR9s
vAbWKbWREzWFm9Yw6XNPX4qKppM7rkHsmSXe9Uyq3M3XwAHZJqWCAedCPxZKvKLS
bsNWXopD2TZC83G1ZhWp1ngtMvgyPZeEjvX0RFQMcbgm1LSJZ1TsfqzTlFl98MlH
S6KnXtvMx/Pdj5PaIbUjYB9PgnCff0PF42K8y6v9czhbwPS6BCsE9v3Kx6EORlck
hcJrRgJcAs3LWTRypSFgck5mlUVTEuBcHnjf6niUD6cNDHZ2v4a22t8/wUjSsjFx
iBsEPP9TCb48NIlLMLeRhXl5hizTGNFto+vhcS25ccJRKVH8di4EZJJT4ywj7/Bi
z65+0CCzei2ACfS+66AIehBfTHGa2FZS6rly2erV120dQHn2X5kBajTR3HDk5YsR
193VY5bDscc1uvtVmnaixeM/+GuavJID26U6r6IO6rvn8khNliULBf0w0QDPDuhI
NHuEKSw1IdwRhJRfvfoW5WGW+bZUP9tWnN5ixPfWvkEr0wwND/sE2KiBcgWPFJZX
QpYwCbe9gjr4Zm0VaxlnN9WpfmUv3KLp9KmV60TI/QiAPm6eEbbN/s7/YTCh27pF
cNONXx3nFi3ePAuEsVxQVO3zeWOsB2r5Zvp3TmeOGvHM6BHu1AjLXzyOlRawULQD
iCKBNswuwO2eeWlpcMh3dRdVAie077mOaCQQkOw9sLKpv2bHKOH6aThBdAcy+Uzn
/5TkKBHHlYJMETT6FRt8jFMSz/pou1sm8ZTDfNDOod2eYhN4ndIuxiAhwKJCvvLy
1ESxk0GrtoFfmngiSpAgAkgeIjJQ64E7yrSvReZjuBlIZcM+zjzdHYZFi7Lr68+p
rsSjy88hljqQ18oLOa07vUVQBy0MaU16NoZ3e9BbMZvykaTEsVdIMFk8UgC9rI8R
+nrKlR7Vt2odKvo0lO4wfMreoGVv2yosk5tczqzhxdL6yC9Rx8+KV6Ojnnuh15b1
OcCuciJOb3Ih+RpRrF3qokUTimsudlLWYxJRaQTf0cDrSN/lX0yV/pzFs+QKQi3C
Nq7q8bMxOrBSXnXBRlOC5ax2arGNHkE7rPS4lw3nQV6U3gk8mclViG8KJhI8o8aV
XhM18Nc82weY7VLCAxWh3+xHGOnqNtKaJhE2GG2mMNzK6EouMmzmhQ35WWOrfXJ9
b8ykzpVn4iVZ32LXlzlNPdbW0QUuLF0cXxWiBZD9DJtsInaxWQc4PDaHOCooT2QM
jnE0IdAvjsCSY0lAgi6/kzmWt1T2LUgR8UNRvvaD3sFLrGu7OGPcCBP9TrV4fWMR
oF/1ARMQcBT1mSG2g1Aaf2p3uT9sg8iWgVgSV0dENB6Ty2HOhL+QMXWnxbgswcUS
rnkvDj+ADKYHPYV/Q57Xrcv927dpp58V+/78Lwho0HM9jpPhFCz4inODpZONK82u
pvZfWOJHDA8bxb1uCbr3sEGvh+f+y6Z3kTF7rgGTmvdwiRvCd4CEHl9GxZ+57Syr
GmFDSGlV9p2frOE1jUqO6M/DSo2iedRXzIAAKKdw9u/1hIMCYqHlLvmKbZ1a4BI6
cDbW4xoMB2gJXb7fctlgu65jCZbseUsJHZlVavvuvKnuBtpsKTWld+QLncN3OO+i
WVjCjDKtewJsQFcD++GLKdMj9ArPl9b0Xt0WI+ztKww1fX3NQpbwdp7v2h9CM58q
Og+Mjch0Y+jnWrW3ac5IvyKkS7dp7tQ3e4BZrERoBSx70IfaBLxjipjSZH5jQP8u
usrUzsD5oHCfF+9ibhJWVxqqdrkidl8ixXRA2EnCBmABGlUDq8FoTSi2TLEGXhDX
GOkNqjxhDmUJpQF2/Xv3Er2YdWuWnXytMCkmuFvakOmTxGJ+zHuAJlxfpaq3ntQ9
8Lc8TINLt7LeQFUMx8H924uQv4pFQxvnrRtPVxkww8I0WR6bWPo+YAiU+h0kybKj
Dqh5nBMStGR4BecEzeGwpwsdmjW4ysx4nE2GOR29qW4iye+5TNY/KYfdpFg6VbJY
jlXS8ds8pxQQ/xYHaAiUGs02VSOHAjQAa0l+mEU3nn1Jq/ArtPGkOWWoY12m38d/
QpsmICHSTIX9KTUdLcOPpgUa7T4cB2JXHriKgR8l8nf2N5WSJ+sDVUUKhm4Crfkn
CgKqcfdnsNmThD1Foe+PtANtpPEjanHu9m/wHg8NeOHYAn7d7fIbbO6NAwTKiAwU
zHhpCVMigwzYxQWTHTCIv7E0kkVSx4WFTzmJhs/LvlzkMsyoAKhns84UcRhZjgfb
tueJ0WDQtH9RfE+I3r210evZ/ONUssN79te3rQCRAVOvdlGGQC3ZqyIHgafrttED
KeRgZkeD++a8MX1eYjsIW/UmwpWQQNIIBwf18kR+1pJQwtG59Hu1vwK6C0l8TlDw
36RT/zSr5+zLmECMnpXuSiB+B58mBZCn2XcZreCisd9J3wwDNLDRUeUNYpIuSbqE
krbyidh9zcVAQ47wFGmSWsqMLIOgGxi3vzktr9UBZWhcJJIhhC+Fjx6Gnc6pyuMN
GzxselqIwz3rXy4LhfbRREvcTqbSmrWiYrtOhCJiSxLYt99p+osu16NlfaBPae+u
s5geXUz+yEgd5rXkEfy6YZKZOA3h3VhNNYuhon643MjegaHNMeZBkeF2a23nofud
nK4lSHh0JKO9Oa0teMH1akw6KDmUWF6i372+sgxFdRokCyXvkgLKZ9sLn6rFRMbg
6+pVAGLK23gefq5Evw9LsQ/KuRGGId3TsjWcrys8cAt1KqxYJWlNaBSki6LlmCuw
338BDcEXFzQugjgfIZNGMDNhNyNWy+tbYJSlmwG/ZKzz3dJYf0wy5PD14Fn7w1KP
1oDR4sbOpNB3Tyl7eUh/YK5PP/g3xgY5aoAHKZDHTw3/VHp2CO7FYt87595hkvk0
WMAUFgEq/gsgfS8rBDmUAmUA/YPk5KambjLEgiJFD62k9QzagJoI0f7buGIFhR2M
R2KAl+MAOBpUQhvrrtwsL9hj8O7hpGcAt/i/itGFYD7HbVnYxbn2z9PNRJkPT9wo
Oq3bIwjh5usDtfZZ9DzwVFl7huOwTZj0xSsDL1esQOlClEJI6OwGGXBTjFHTtn4O
Mdl8j9kgSNsbs1aaIUeeH7Dj9ioIOFbvH/2z2QdYDmXPaaZRCE5KahX/bBnX4tdC
dTj/sWnLuMVPUfYmKN31UzLROywJA//QFk9qxJ3BThNPKtdYlWQ8O5PNjDlwKx9/
Y3zLyh2fjRbNSy/xZOENRmFhuysz+cpUUklAtFoxI2fS8FH6iqYnqeZkF2TZgCOL
CEkdSSNx2dAEdyQU5B9flGUtSWOsCSZ/Mx6LtOR1MZvwb82pMnr/nv3pk7/N85Xz
bJW4puUpGxyKZd1CfSDPEkK7RuqucceK8lug/g/kpJg6CZY4aGzQY81qmRRQjvu8
t3UZyTGwJ8a3NUlc81MiroTF9EpqKDUJyPsh6oX3mrjpI+DqTlo5oE9vMBk+VuRJ
YfNfMBnotL6855XxR//AA4NuztdPnPtTs8HAMCaY284keHp9u7aTP+kEtzI3b2Vk
G2awXOaZTEoZjMi2bGof8CA0Tm5dDRZMd66rnd+pP36Mk+Tm0p6d5LaSx+ltw/UY
9bOMTVZd4rNuIX/4Kk5KZdsE4GawbweOmGcZyZKaIvhOdCL9B4BdlIptX09wIQnp
kFWlBYwXmJbmmAduRSHGdH2kWtqotV5YcSMOpezX1R22VXNdsFEKtAJve1mGx0Od
ZOGV+kc4vUdtSRDlE6wNhnrGnnJ7OpfaZMXkUjV6/bWI2c3XCUdfWw6PILNbcT+b
oDkFjJW1sWuDH6SSMGyJhYmrdNQxciBSyWD6weSp/bbdOTc5QRv1eFKqflolrKFH
arxC8Y+SI2rxsjgS5DsTntl4vF6k4wXIExfbnYtkXUVQfQGveqaI+btVsSSQrYFS
8U5Yy6ASvKESUcOWUIjWW2ouu+kwZwEEs+4prPH1prMIfmEKWJFpnOjtGx9+XQOx
maplOyU9U7+PC36XVJJuYWrUoUr5vU6Et+fcvhnGHkbzHy8oJCWYp6KycvvnhwKq
RhXoISpT8tNTjj+bjKaCUlsvgN7ZJIk+zhEUmsY5tfl/QBkp2AKhvIEePpDlhftX
o4+0Xu/LNDiGoYXXU4EpcgNJtenKaZXLrBai/GKkEZBhfq6xabYiPZaxp7EGczKe
yxvu792YSuiyPjXySZPaWEgITK44ILc1CMD2kxyi/S/MrOPOlDF/Qe6zJ4YrewIR
XLtikWE1HLT5GYwFWgIzKOJGpmCgQVyatBWlX4CIe+NMjIkCjdEGGlreh8uvC6Wu
CQVE7xGbbEeaoJl8fh/MWlwc6kY99B/T65DIrJmVP9r6+/Lrq/WrY22La19QL/W4
5MF+6pXS6lubPa4IYXgCLcAn4kSq9vu/knNfR3n5FZacRFndEVMngpMUsmZaWsD6
Y7X9N5j+Y7eKHFAHjMNbq9QXaCRw2P7hiQI3Mm5WNYVLzl2MIhzuHcPlfhD4pfp9
MR9AnLklcGid+qsbLu9jyoOuQ/UjYg9tYoFfjk67iOmmjIdvkary82TRW3E5cpSj
jyBJbfFdlbeHK4fhHgrNPt3j3H9RFUWYwme1f2dreiHbjn9QTBwH2M8CO426wj9Y
rIs3TspkdpvB6pwnccceEgST7zH3tXTWEm3LwVWzq7oCALjE9eZ/vQ621CxvfMAf
VkOrOpJ6XBESEq5tx1KosZTRknorpRaLscbzS+DITbxYslL9HdZMWoe9SvdDthUM
3zpNExWCIRUnr7KhhNFLe+gBhuGU/pM8OTAmXCcFpUWG06PLhXxwLM+NzC42qTLg
0ZFU9avMJoX8WGTqLBwXOlw9sdEdkGYmhA/shJSarhtdqncFr/7XDzuzlko3BL4h
DCTsN1SgbN1JMUCgjVO4dXe+EDfNgleUypmrT8BTTBqEdUFbRbgFCHLnuF5QRfH8
s3BsbYZS3M01n9qpV74gL88TQa5ChaxC4t/c8vYH/VBGJUIOy6JVySOcAmkF2wAq
DlDHrC4KmxwxQIdtdJX+VKkiMAx37WyoXbxX1UboSPCDaCCps6nxnZbVMwk3fiZS
ONLZ6RxGqm/6iscDyD7rjjavR8JCZpRXXrBuh1eN4E7q9yZFdG04hT4WllXpuwTe
5/YIxWfxbHbeELiTivdkkOZYlBcH0KDwjxUqaynNqqsy/0wjdAE9BhvIbesWXQBY
iAj/XnVmHiRZI2WjfDvfG8SY3l9oDGOHkmD11FTQdk3LqTeXu7L76q1gaS+LPJup
ljTLyhvGUiMPmdJp+lTLdEnE3HKHBcyf6HdjiQJUs7c8CyvSqRcfdS3B9HePMy+D
Hh8z/CA1HEX7X77UEStMxymd7qzC0fV13w1V2zDR3UwM5rJjns7V8QUmofod981X
OSwCbER6qk+tfZEYXiNVGi/Ifcd7D71DpgcVPDCbVa1vG9YrjEsOpegjRBRKKoA5
398ChgGg7jJPUYe6cF65DzpOG0HF29YdudpE89nXr/E5NGYWvKGSlLubPT/6Kcs5
v8tucVb7gOCyjNjc+e6DnBOQ5y6wwUctPqYcX1eIl4JijUukEn1XhOafrmCNS+7v
pexBUlKFvD2fvguC+X/DRBfbLWZivyvRSkT85DClrcgCQHC20N93P+KwfRTF8LEw
MtJSwi69CHD4/+KfOwu+VA4oTAr3KeGP0iIh8c57lwmva/mpOthhtAoT0nbhK5SL
0BkqP4YnHMP7Zyq+mDsOzZb27Tk13YkRPBnEvcBVmz5uRQfjkRdwk8IyzmkaT22n
2sKzcoA13yjHXHEQcFTeg4/eEgV32J+2CsYqiffF/ShLV6FuDBmOsIFjj4VKQ93g
iu53XN6BVWIKsFZ8PdaWFYonI8/MoqQ2o0YvW5zWrW+OcJ7FJSMAs1Tglse2wzdP
Bvmf0vTvqav0QC7fPQ4mCZTEPkSkOFcv10LqPLUv8JZDxcB0V+2K+kkm0N4hc66Y
JhtMMahC4mnKFO3xXd5kCLbHnnIpJX+AKsDHuRhRFfpr2uBXgIH9UuXPYNM3DNNI
v4CDnLBZqMHhaYSk8JU9+o4UVIBsI/KQy5UI9n7PxZaCyFw0djPeh0CobNrRehvF
PdR8Zrv0XA3/nReYVlSXew/48rvNYS1XcEjO6iVlNhekf7qvTorxeUavqsRfssUc
KxGyN2cA9rc0S21Kdq6pJCPFCa4NiUF5eH9kecohTWRP5fxJJheLLsHqxCHP7SDd
pr9sMU1qnFDD2uD/Zpqk0KnNnsc9Rqnop6cQl4Q7SCw+FJjhOY059lLt3hFtdXjv
EBFlXVzneAt1xwAd7mYE48zK/QbzWQQ3EdKVCx+PnHTibRDhn1O8AV/7yKc0544J
+Q5ogmGCirUifZ5o5Vf9s8VTAhq9acKFBmZnV4L/Fu+FiOnUuxiFbeh8L+j0e08T
ElGBDL6n5AgcBx/uCZCFiJF5pZ6LV3kpnPTftB8KH0qdTMpoO1szUa+waEZWYIl5
580LFC9w3uvnPwoMlK5546R74A0BVJ/1cHzoUQWrO7OM8JPLSXvP0lM8luyPL09B
mUBje4LhxUPIG+oOVvvplQqfCTfEisOwEki5ExB7fBsCdPktpL1JmKpbGZJo9IAa
wlsLsqH1OrL2fPbW6O6ynxy5wOcjLa1p3mjfmLol9sosIG/+grie/wyqW612jdWP
ezu5zFXzm7PTqxjp5GnYfc3bgJZJaXidauJPqvVTECO5CjpvmvnIYG+N5rluwc67
0U6rxHDGmP22Mxa1tQ0Yn01al4ITnN4tjg3oCAnWEkbAyA457LEV0xYszywFYpKh
9+bmXSzB496vbYLk31Ln+6K4K33PRBU8BEdwr5GTrZtiG9+dyTSBjHl2hOodUQqq
4bjwI4CQflaAx/i1iAfm08W+kfgZKOj18Wjm/JzHN/tGgZyUx2cAk++CgrxljgWF
4lupRfOKMP3Q4ILKOY0hsvBe4KPynL8culNLnm3ANV93KTu0hs63p2dV66g1f85k
QR6+knvMjW0zPlqjMiMI7Bf5zrQje9KIpMRRU7wyQjQmhrVNpx2WO0Vj6S26eWjZ
bhoZBDu2EC/gCzF/5Y9xqipAKF/tino3FYkOwUaJUZnY7x8z9lGH0qpffOwt7VK8
hWaE7Fvrgk1NAw8pghbcbdSSSQiUoDIGze05zGxNTRvIbEvZdP2lvdVL1OEBkNt2
ee66aDq2mz13I1KRl85c0QRxWzPhnMLmsJuyyjs3o1XaSV4WEBJsP7OujFDRKDV8
DU2QO7Rf3kYET6BISkwOF0HUMI6tW9FguejLo6WlNCPD8bwotAUVE01cRaZuusuR
5hK+J0xcd/+/ShAtlQ3McxHywzMWru2iLf8z6jn4oguAGUBeHCUruwLCWMDgZQM6
AeEmqHPU4/+sYCtC6ShYNqtuzjrjaEMzxInCzru5/LWUtt4zSkjpNsd5OcRw7QB7
ffjaJ5UxwZiPKDzRkmBLwW6FAYVb5wRSOeQ6PGziEYnrmiuzYG9WHwBgEy/Z90ic
Cjqtx1AOOvKnj90HG92K0WmuvT1L6Lt//o83QGuPrt1lWkZKSS8b6L3WQhE7ki1+
QlfxWnctut+l172eEYKH56KXcbAbtYj4KJo3m5LeG7dzEs9j0cU+2WtgnkKwBgo0
X2CvWqVVh0JkGsM1jkUTwEe7UVsjtmahGy8sHbfeKrxaUOc5B5frSfYL7acGCCPo
FCkQxJXA01N3f5Ot8FJ9i8LRxLi8sKp4x/Ja9flW4HHlZQUtSbrJhfmAHnOolooF
8Ys1p2Wq3XItQAIFTUsekm/EPcJaDEUH3Tk8D5Q/y6k9HuBLwAxd5Dtc0YmhMq+i
TYBnhaWjh4dXA0xpR9xOkxEtTogTATYO/ZnAIMYM2emrPTT95tFjHV1vl29+7FRi
h39TCSuWp54UwZS9yfjxlKwCRZEsplI7tN216BQB0eu5N3ho9G89tJq3szNTZkks
S26fWUIesTCg6jz6imZFnCQ0vXhmiql3/dQZ06RLDAAqukObutsD0OrQnvzKx2tg
+TFAfi1cvNMv0/oRRd2ip7r2lZ7R40OmkaBk98bfXeT9WoH5hT+0RnGauPgzrDrt
x2y2p1gn+DchKOpZ7zwFoRS3gmpRpjfuMNhnN428LHYn+2LHSy3n5mxiL8RB3Xw0
TBrDR5In7ofFC+/eXkX/uUMucY9sBwPoHblXdzj0Mp/Eh0yOAwpLvj5YjlEdWfqa
H6V7knIitwO+stEm8D1GrMqPzDf0g2Wp7IxbYLuwWq5SrjRLsrwjZk6eFp9sJXJE
/hOLNRNn3pipQaK7HaGOLh+EqpxOWshfHOObtxkm7JPSepFFni9RV7S99/bbdUnF
nwXRE8DEcRz6U6UDkqD2G04Hsi6MWzku+VsNuRw1ahUlypTTaOgC5g4OQGnSLYZ+
q51VuocXyB0YJMmVfbF+L992PHpHbhrWcJCviCcHRUIiPbURU5vnDIu7Ypo3o99z
Cc/DlRHb1fqaCDJO662MFTmm53zmRsoPOdrYHtZyRkIKfowZ68horRsFOHTSXxqD
hGQk4S0rgK8JaYG5Fpg9g4/XFOiD/ib/1kGUAv4U4Uu3hNMmps3yeDv1J2D5vyr4
44paCLkCm9eO4rpq+OxnEyg7+53U0jwVu28h7nIm+E8cqJCMBaIATfqZXIdU/0oQ
RU2xbEFWsnNDhqrOSKXa9uI31fWx/gt+ktCEiOiXBGMwxfwP8p3cvK3giusoPUnB
XvL/Ddmnu3k8izrq7tclqmhBib0eIondknacyaW7SnWnn5XyacUZ02WvAwgDRg92
KYKYcaRHCX2M4yVnFIb9mitmblocAe7kW/KlpUGgmynhQJm2qtV2IW+7hTi59BcI
FmRmJr1B0xIhRzi/JqncEH5DzalZdKOKZdb11bh0DHaE2NQGbkYjxPuFCQHGtD2H
cE3I3J7PkSvEBr+6xeQYIdappETj6MG+sixCeDeVs3QV88If4F7U1/t2TOprNypK
6x0AoQGjzRBvP7+j7lMb6JH+pa6pS/9SmPYaRY/feCY5QWvK05B48qQ02IdO31M/
JxQl3PHaPdhIOZzhiWYeu3wPbMiG/xfxqHwZpXMgtxU6u9PJHHOvrf5JUR5NHUou
QIhgGAyyk+rjm737ueeyk3ZZqrs7iStj0jtTuVTFGpi3oznNWSz9ux/4XTuGdUPI
YkfZn57eEttvPYy9gIJtf/xV0CsAF7WQsA9VCYZ7Pw3XaSmWeG7MSdMfehWLxsXy
LkCXlsg9BqPBUW3r+KxrfjlV3+wgkNfxK5JaMSZXoHAFyaZohjt2re/K1ejVutHN
JcmTJ5kAkc4Aobbe/XPs8IFxeLWf3G1l9XX1oD+Xvd0IvGn5x9m2lImhb7dosPET
wVp571lJAa+mjQ4Sv21p9eiBSzFDxj/CGsfpYnobokZinOP3lRFxR/nBvsPHaXiQ
PhJFJR8rLNLrf5GwgdfP/LGW1GNaoX6uLq+W7zGkdL/Wjr46knL88fayGkgcD1T0
iWUJEkjHe3LmdsvKID5yHdMzBhDWUiSlA4/875ZXkHYWxjKIuhsvoco1184hdbiI
LOomdGutBRjgHkIIR5KRONTPN6pRT64e5mvexnqDfiX0elSQ9pu+Ito72vbfRh3z
mEUsYkYWTicht8oWO01M40bZ8wcpx9cMj+Yp6ezfhNQGxYz72AR0RF3ckgsNvc78
Wmdn120mEh7Yf6k+eqvzIhNt1hN8+qPVt7FI/jbGANvNr5BH27pStmzS6r4JHplX
NjtAooejs5Jy88527hg08Tnitptwd22z1tq3EcQwTRYKrNgEtaozC2hIhchFfOkV
4MnWDepm5QRBuJ9SLqWj3ZwiVJoNh9NvvJ0qD61kKsQU9i+GUyPzxoYauNrcu8mf
ijYw9jcbGttJcVIsWBviaWvENwx5BLNS7BDc+P8J+qE+uZmyXfQVEBIUogcYTKkz
zqz/ox1XrGjfYVwX7AFb3VPC0/ALsP1s6fcuwaM0njHd9YecQq6XJPi4Z4+eu1+M
hRIifrmVk4grM2lAjTcL6pmjnQ3J5oGcij795oSupXcYBLyXsxGmo1edulmXZN2A
MYCaVXAIVJ+NMQGhtNy6lnjVANnYPLvN/h9q8sm7i3qcrByV6uDJmn2am0ONiOwY
NHiLhMUIMlG0Q69gkdhHfV+1rxHZKCQVaXEbTmS4BPdy5Zi2ZlnDAz/lErNGbX2r
oaGt+9s45HwzKUKHLB3OLrWlQHbkb9g//hDQQjhiAQsh5/NuoooZ0gJtIIXQ2L+m
AzowVLeudMx5D9TApOjcGY4QGtiRZZ5J8lSmItsf6cGz9xn+rvcbH+nzTRjoFX/a
e8MBP1571Emi1r4f7MwJzm1L5dTYmu6QRDlPBFJSS31K1nzb4mM70spEQnpPF5VF
j6rvzcwcGaHQ1plMT8iSt3s79L+MVNhQpJ+CJLhA03eX/ASkirV8BYEdzCD9xkn4
LJIqpQRp0BWyh5m6ly4a4HECSB+BATXp/cGnmJQo21+GPkMAhl3XEHiD7S0+V+7/
FI0tO6KMgY4BMcYGcNDJ9JkIzFDF4vjxR+UK4SmY/i8Z2KRRXwK9E1j2jn15HKSR
/NIU7i7Gu96hp4y6uAWbG/zhLF49f7WqwM9SZPn9fY4jsK9gt3QyBXnxS+hs+AjC
d4WUNbYx5dF34Q7+3jU846YPGTa8vyYgOA6taMl2IF/cOTOS/BeG+PcukXLcwNSG
xI3GKPcLnNYeHCyBysrLWHbooOhcpO9cZcqhovZ8PZp3+QPA5dn/UYYxbf9zQJPM
oxMg788SyMFJKCfIaS0AieCjsGS5pDmJ1l9TuzQ0Y+8sKsi2dlCLDVbX8oNaapBx
GJuwUidyIHeky0fMx+60KsIe4WqdHQj8Ke2PKHZUh/VqFbLwAOZrU6XzpOi3X+jr
7yE4SPsrYM6/DX8yNc8qhUqRDMPhyrJLHoUTuYgre7LefOsfL4OnTuhwZGmhYaB0
f28Cc1/AIhlH3OH0MVl48XF1NCOGTrwlos87gFc4kH3wcGlcRpbAOoooystRS0Qe
xGM/IndrL65YNvSJEPexozryr8/mLGPO4pgL2Ujj5fu+wibHArf8SKM9gKr6X/JS
PDlNEDFH+4Uud9YGVtcIlXplTy2/MV2+fTw7aIN+whmusJ0UlllOEIhs9DN3S4ur
4L6U3yCd+9f3nbP2Rl7vYKb2mZDVYsMaXMPdA7WCiTgD84vFNueAPe+yMdQuivSR
lhpFzM4Nr6asCKFOa23cHJi/p4WVFYJIhgLD5x7qAsdeTpsvuEkwFygIsfx9X11q
x//iQsMa65RCZu7XAmoQz9sZm6cvsKPZ83EiwOarhmJ4U+ZYkdRecw32nLWix6bR
lP6F9ZcKqlA636lJBZg6WwDp8HtJIwQk/uf6F9Jvg5cxIbAysvCJcoMbL9+JNhI+
SBfFcMxLq/2IkC4/K+2O/QoAUWZmhZ7XP1gLoyM6Hd4PR4giSPh6QQeCou8BV7QY
IP/+lTJDqc8G5yr5Q+xXQnrNXAVSnFGrCPdx3qOhuN7XHaBIXV4JOYiq9r2Kydya
OHkYhqfgVz/sGJ5ohalaaNV3w4GnHPfrYIl3RFDRXNHMVibivK3ZJhAkOh2ObLLt
UUSESS+H0RXlqEf2cyNaSqEECTw15/RLBl0h9dOGXewF5z8iiqyhsTnurAMajnuM
AdRMGKgH8Nc/54KfNNYkxDrK1L+uM4Pvp11BjDf6Vy0C9P+EIBKECVbkZG6+trGJ
cBtiZpxbR9S6NwzNGqrHdXxuZalMv0KoUqsMDWI8UZW8cvwq8rZyKsDX45cJdlAZ
v8m3qNlMz5+9CMvIxkJtVot7p03COAh0EpUUqxVJoQIK9XBfXyVthoD8gXz3Yeo/
Mbdd8YfAPcOZDchLqYxsdwgpBN3MGbpSYPe345oYFcPG0890H6QSmfwQWzldBO4x
o9hM2W00VIJw/am04yljIorBP9PXI8yECYgvA2y5ZuT4mUGC6fRloMSJvY1ojUu3
vyK9luarAOEqo0H7J7uVir14pR1YC9WEx3FrvD4PqH9oaB8pGWFeYWngZeHDkO/N
sX4+XOO7islAXyMzIT0Rfn0rD6HTIZA/kVb35jQTMMNQbd2s51BEiN114NtZCJ6S
uki2Ko+2Ipq+SGCqOVqck+lhfH6FrLtnnkaUDR7DJ2jt9gxoqRVhVejFIvXZ43I6
0SVgh223NHMULeUgb+KsNP/rksx//6icf2EUW4abrYAh0GZbj1XXSipVUh/6K+PQ
rBGP7/3779usitaM0m9x23UUJ8Tn2QAyUHLwXV4wFo0ARYgZoHulPB+ithtoCB4o
Kv8Fnhghfy62TXUahe14nDl0lZVQ4bekb4i4KTid/fJMbvc/Kw/QHfe+z1+mFBdV
Or5HCIsUk2d+D9ZMbzGUGzcEiRwmq+f7+hr5vqoBDJUIuQqy2VaQGAzL0V6U89es
N5mx+7efvrBpNDzlHFWdwPiLpmvmrwXeylTSTYH3Ptu6sI5NdZ7q1cM/8pXpwT5e
A3tczViIDoo8lyqHMg5nphOeZ0IktlJydyNPcg6V7Prxr/ACZrasvxms5uh1tECj
yhrh6yb3umw1GQNVpb/Zd/N43cTOIQGoYYF2ktmyNo7my4kdwzbtNNJRWT6eRXAu
ZoQhp7/Ex9dtT7Q/1FinKMox8685UcIrp4Xq8XYdnaH09Y9ymFsP/hmbf/9LOzfZ
tFd8MVfSIgfUQibMRj+uWzXFTmYGmlj7aIctKKUDTisc/u4Rl542v3HReNX4+RpW
kZ+w1sPnelXMk9raingz3LYAxqQl8MQbdSwAPcCn2XznmzyKdPZ3uQ+JEdPTOPiJ
SWFkOCYYrkQxyfNBvAcI+DOCHrwEPsbHtqDqlF8bar8WQCAknlAZbSnju27LYmt8
/YG6L/msMbebnVfjI7wq6M7tDFigpipkaf11dbMbbYxMmnN5TuUC1wLYAiCUnzUG
Rxyl3MM5x2PLgi99Pe4xzTt61D7sz+Nua5xEjutLRpsgv5rIvNgnNtX5wTie/LqL
+fxsmNg8BEyj/ARJKqtzdv8piWBJ02p4uapu4tAbUbj9P06OeqmZ8nlSGvIn2wVR
l+HcZ8Lk4j8BzciwC/gNKtpfMQiD1lC8yGYjJzyHL2qIGcaFjYdXytss52Z5+h13
6VkCKrZo9KjRv0/5KGR8CkjslayTQ+mwBCcLGBE+bE6u1ws9uLqZetoK5QgNntwg
rrO7IBPId0NZj7Frzbn0rss2aDGbEhe5sYore+C5whp5ydmtlLJpCw7Yx3M2CSgi
6ndZe2eWAB1icibCW2kvUbU2lGRQ+3U+ZTXZvs0XCNFI9oBKLoQQlZF+nfinPNB+
LI+TDmwJgd5fBzRp4BJc+NjGYefYBoZaKixRBiOUbOwDfl94tQ5mNn9mqU1W5Omt
nyx463lRNC3uI4EiPn6LvcDYeqvQAKUbEBlytpOUPbuPnx8vmf7czVpSke1D3XwF
05/5ZHjQxHq98vtkTQ9uDHP/0HGJCSSJx3L7eqwc32yHyh97QMY3Mxrz9U/nOGsa
h44WD852ZVZ1fuF4Q9yYp05OPFJmi/HQQPbFYt3O6u4AoI/pSHWy+TpHpj4sNuKH
9DQ/SkGU7h4RHbAM5Y3QOpxB4wiP1epT0gy6TMi9OUCf3+k4fCi/hV2VDvzfk/oH
pJWp4ZAC5iuVsIjOG+7kKWMiVJrIU+xvEFEzTDNqjgsGGzrdiIaaFX2z3BkW8Thq
99Tz6FSeSDcw3KxHqXnoVA+1GhXGgmyCftM6HJRsdqFvqiFeJxdDt+v0vSodfLCv
afB49jHEs+mP+dIDgSgryAiGpQJEya7U3cXb0/NVoPrDK1sgkt+nAg0SJ2SBVPkj
PGD5Z8SOWmFA9HiWnrM/rTaj5MAfCMYgnl5aVnQMO/6gGrGFdAO84UfNyBacNCBU
9BlSTLD2iuoh9M2YwTl4SWm5dUuoOpWqYGMHXJvGhV/50/X5DP3xBBCP2iODhosH
B6MLEViFxWJXtjRE4aZ9NEEQd4zwHuikOLd4K4Q4AMLj7YbF6G9cXAZ72r3maqqC
xmGI9z6M5jGNsfEpSivG4tBL2pg5G5HmKLUhFRpiYTZnMmpT64mb/D5J8qnZW2EH
WQxn+lyaJGGGBGWZDem/7am8dpmf6x3NgA/+dxHgP3bHL9okEYLy1AjV3JxFvlKw
z/rx+RcCtDDXuHz4tcfsKEGNaut6ZdAd1vpx1Gz+8dXRIXEd0sLTc0dtYIqM7+aP
5uDH6kote2+8CUauXbq/0R/1xYrVe+G+YfDDtU3d4YsVov/G0tdX67hsRf5VWV2o
/9uflNamzeKt82GN39YMGBtVtZ8Dnwp+OWGhqYFi1wcJ+Cy79wL3TO5Xm+V7VI6M
JzsqpYRZRMQvkztCouiM+y5wPFoei8NtbocBEH28lPi3/gnsWpOZLo0aRo0QSet1
x1ZwWfbaroypYgmIR+SNzLb7hWi2eil4OiF3CxtX7G4ntMhFw95CCbbY3x6raUoW
LPVdkCnucmAvgB8XH9uHxA+9CH4d4x2G9j0gEj2aAxHIRz4sOZI/8I9dRLoR0b9J
EPqhOyD9okvHuKQxTbq00yZazRSc/B9Gh9EMMnDsxQ2zErBr9tuOR4YA8vnQwiUv
vqrhypdIsaaFN135Uks7XLUpb4gU1rcwp66XYsZ4RDNS9wpUIPVebgq/OtupPP1e
y+71TWY15kf/Ys+ayqI4S7OLE0dpeGa+n4YU8+pgN1QdCVZsjy79cBkQEK/0iGjw
Vjz8RwqfR714LvmzvIAuTzIw5iY7+C7cu20RVrbZ9xVsfFD+lzR/todrWGLQ7dAH
3BZGMU/OMKicwcRdsf0C5+BS/mMUIpH7/lXttMhhX8lNoBCrH0x4/98VSXwlc0RK
26pQjKDWVVKHGnlZ0/Z5F+2uWRoaQcODZPXQ/1QSB9kB1Eax7oLe2YStboikDb3d
DrEmLeBjyKTbl4lVKGjOZfo0S0MpkWH1ttBmfcjzzNHtL7lrgpS7TNV3a1rGR+Qh
S192VJTbmphKvTZPn6YSl2pJiA9R9iPYl9JHW9wRNcZm6WoXGeIKLmNGL0FsN8QT
pxHOn3UO4AoFHgRKUQCsQlH24aAA9h9jjfJmtVlVt0dLZ1feHcmMznFSZhlZXiBT
XGeS9Ke1xb+omZmv3mzZ1fm8tUeddV2HKMuzv+u7i45e+HmRh7ikHUn30D/hiGVr
iQBC6OcmZDBhU2FfYNHsk1KjUzLAhsluQLoS0NvhOub60IBlQKsTipg40Uuslk2t
+cuGYSCIOX1NfgcXDQ09CR+Sz9B563zjBwPTsXd1xjQFU65ZF51ManuZB6PD+PLf
l5Knfp9tNDvXpqsc2knKpKkVLsVZyGH/ODUW/paqEsmLeoy3gG1nptlMv9T3tsXz
MCeMrsbHQSl3feJ5Uajs5TZEwSSmYB9Qc0qOk/+E0afmG0iAbXC0Pl/2voUmlcQG
xqSGJUTyS93T5w0aQnvt8GQTNUqvR/oZWfyKgNSzMbKaxb3YCVsdWAMeDoTL1Dri
4IylIEdbVqGylSc4ZBvAIyT//V0oIMqTI/g5L6TE0m/AmUOu7G/2+czhs+ubfD+C
MPTt/Yf79jbrsWJcVglHxlzNRAVQQWODHlDYyidNGPtb0t9DKHZC3Xjwh9v72QcE
dT8QZlkNbEgJ/SsWFYzT5e3MKrs1FZjCT+RIu7uPEAXMArjGfL6uZtg7BX34iWoq
nPl7wrdA/LW5M07UvW7WnH+I29/3SowFOk8dkDHqaWTDyqlHeggI7i0bzeHWux9f
BF+4SB/Z2waLIeNs9UBkmWCHSPWoP4EF/8DnQHaLKJA638RCA+fCP2L5Lcww6tAe
T5rl0BqEF5Q4iP5Sz/6o44kMIlbVT5NA95eTsAh2Hf8gNxexWo2uRM+XkRVNo/k6
YjfZfkA7s3ggMlL+9oVwj4BbZ6D4Hvnl4LUBAG8jDjWQLAqYsZAbOVOajSp620Gs
/kgkIrdHwwO3HFmoHfsNzS0irBmwyqXD2Dz78IoVMaZP7VF2uH5k9vNgwZ9fqt2B
NG/WbjT7we6xuVNts7TOMQ4AVmYEx6o8GIw940mZIH5AmmUKioUWoSKKEExRFzGK
9Xgac6uutcr0qY407v1ZeXx3Vl1NTe3fzBCHQ2/mg3SuBNGPlgcchs6FcRCkEGU3
SgeocVUx3lm74Q6OGV9kuBkMDMxAr+De1iW3gpgqtEYB+atpzsVz6cOPC3mb5zM3
crGdxNxPfYQ0J0rn8bPiyyigQji4N5/gGvzAMv3I/xG5fdyAXrwwfbf6vPYkmMMp
V8gJzt6W5/F30bvPTHTv9moTOUdQ1tXS3USTxWjBK7VVtWaD/7yGn58RRo4UFNrc
axIeJ5bwiUnMLwm3/isOInJar+jeI5oGAI7I3GyERnIXZ/DacE21zmWJp/W9hFPG
Enb+IYTVbqx5UW39HwIBJrtRLzqQRyTix3CVqoM7rmv7PGlRCZ7zrCzIZYmgVJlz
5UV+ysVBGMQzt7uciBznhnipiYDp9A63PUWbdZGieCGTPVLQomCoON/klELbnj+J
8FBEDlGho73hXvMrw3gr/+TjlhtTeh79dcZg1G0uykcOkswJTIfADE5yPmOXo1QT
8Wh2zrpUQ4fqowkfB2Z49jswnxFKqkaq6uQ1mlxH/P6VQJSNUFU0Je4nFlgUA7jG
ZGf8H27N5OaYZytuDFJyJuP00Zy0+P1ydF228oNh4lGomPPHPXO8J3E3cUfpctKZ
YQy0a2N/TLDk5LFQ7qEM9ZNrGjnebOiMCyCDODozSUtN7Ttr4cgqyf971geIIai0
3613mmzy+pkABRX76bC+UlxG3zc8owbbD/XhWbHUy2+H/VWmaBcdXnbK61KrVh6g
oMCbWAw7882ZTq8tk/sIsj6zhiIvAbW/2147rmDd1LN65oevGUIMdtgvqFzoZV7t
opi6BCRc79L+ALiOBG35v42LZKbOKPRyh9Qtb/MywpvzO9dpnVwyBaXTQMpIAEPl
mAE8XytPA1BB8ouqGrE+xs13NNHt77qYzoKStDgmM8Uq8XMx8DBCPrJmlfuqZzJk
SgngbaxPZV8evCaFnbBVKlyvrCh9MeHOt/kn/Aa6sshBlQXRZmJyAI3IVQ6egSfm
JuCqib5rK3qP5BxckJ1duJTqTlIQGytYYcBMfFAkMlLVTwqHbRWmrXUrdWiZHV/I
4ISY/A03u0lIs8SyqEE7SCpIJE+kbuhSTEzcsUNaHWIMH3z8x5biTIFcTqm3xfZo
Ddehq/AHBFCTwM4h/O7kZIb4cN3Ae4BSsNJekhGTxnpioPBehvMoc5j03x1FMntk
dkF4Kmo4rCdIK8i18T0Uj7hH1lpbNtqblNCkbYdWBSDUltzFONJ1etNtKcouXK4I
e4Ew8sVgrVHTftnz6VNWek8u0AQMMQsmkIFOnUnKTQR99Pw1cEOqFmEETISJKcHt
c/s1Z4VVdgM3QNaVVNE0S5G0kcFlK/OjXqe5ZhG8DMO6voyTjFj4fY23kLRhcn78
leHjUiJPjoUgl74HUkJ0Vo/5Jmm6LdbstM9R4SqZXqCD9T5I3SwR4ETYXTY4naGI
JFBGIN2/sUrkdASNNlbMxaK/dxpShw2+QWzgJRrwZkk+1NV+EfHbeVzIbnfRzl/5
8aMh1U3sD/uSg0kXCAEg72fegLBhyL8oSwFC1QNu5cBOgI+kEY48BZBwS9CZV2ul
wPuVY8H3NwfEkk68Ue7WOgwcqeEkTO9Nr4CNSG3Kj/4aidtrZzmi2q074af6YfSE
XfMk1FgvAUZ+Xvfiwvi8h5xU9zIGvnf+EX0s26Z/1owPl/h2KphNJfO6gQJi5UnE
HxrZacU1e0ZDnKuvNrudFwJDIRhHms3UVrWoY+OGomFHVwJrVoFaBC5YsvdmVCRb
J0g5t4+aq+eujnTx0FpPEZLDFStKik4t3FvWcHQVGHAvqEdWIWWV5IbaGDs1FCUa
LLcgq9UgJz1BU0RXrz7bXU6skLYUN+0nQZVnoNWZtyGEfs1zf5SbOhB+l+QyLL+V
mFpzAZJrN1643uWNZySLBv87z+Xq3RkUg2Xf02Vod58Lb3gIST4Jy4Car63lKBRf
2AfJ1jAK0dfBT8vS6M8rPNvegDhUFFUIcXsrr/VubStrUxxxIyalg8KbhEymxFRI
SevX/v+y8WZt+wQQ8+BefqbCFCt+t+smdLCq/XgJznzcJuO2IsPBUmqxx5QRr0Q0
x1r14JwAkPOamiZg4jcMs2rUl75y8XO23+sx11tjuFME2P++dIKxwmCamqFegUz8
OVz+X7uq7890wSbUEoSuOYvrYLbvhoihDkZFdDHH4of0KghFTYw4bpZkBkx1/IOJ
7jRZGZKkHrnkb1MLlr1QD92irJd8gasRHXyOVPZ+xul2wUs0pOf2rCAW/qNXtoDO
BVVAjxn37E+aVLDMnZTAQde9qsZiCF6UObwX1CdJmJh1C22xTAQt+gvGumamBbDO
t1xMWN6JMYnAar3gU0ucsJbBp54HyVhudZDPdt/upqWBxhChPyV3gn6vLhDtct2/
CJba8qx/FPu+pCTLo6eCf1eqY7tUdpjXU8KuX78kgl1dQeXLcnAfZLomPRxUjPKU
3L9Y8a+EGVtjLczQ/SAiM0pNfiNYemlBVuOTM77etgpfYvtWGfw0eEmg7muP2E2f
k707n8ViQwTfcMIo5htz5wa46xCZ07c+lOsbDVHWwifB+rUULGhKvNiVvDhLksFY
h9nhHSJUIue/Ki3tKOjT5SmHkqt31NOLtwEPBYqANB2b81SVOTRcPlEEXV14Z4JH
7bRMDFSpaetpEALdPpvY39kZuhM68UnHWanYAO9ydGhqNdEoLghKoXwiWaEV4pE7
eXGt3iIjz6H2IchsBSz9OuEKXDHq0AUnGeUGv/d0mqEeIA9c+IMg1Riz5E+CDrG9
Zzk/z8o0gQRSGtqv7P5H9OSj8YQ0YsUdnRkie91rxo+bA3Zcs/kZ7NWdpK2e+/Al
bq4Hjs4vxPDzuusaIU+iSnL1xJG25kfVN2nWXFppCd1BvKVGydIh8zPrQZL5jWav
ki8+Gd1ntYXEy8mPfulEjO6f5j+GSuOdoi7n8x9tXJ3NtV0PjlLmbv8Yif4+UY2E
Y7yb/wjjHd5I6P2k4tzr04aoOZKz5Ynb/9b8CIsL4rc3XpejOg8dDG3aAdlBWQqa
AfUEToey1XhygYc98muiE58YODNRzqqtqq0b/9YcqUHPIcj8Ty23iTUpyPTGnfGO
vchKBoq4Lasz/EKNYVDdZ7OIKKtGivkpnJmlrGSrP1g/zf8w66Iq/M2HJNzXLzvs
gPH4y1SVA23ulW2eF1cqdIaPEJrEwc97nLbaywGKOx1XREWmorjh8dkmCpiSvtfS
tu9j3BVWyAXTzeQ9+sdf05FQoMsRXXQAa0jNfcgP9K9JX88tXKUXtQV8P9PcibR0
WfFSacJHvdPsJgxfI6LUOIDTghcMUni+Blpf7mE/MiLP0PzlKyFSks0xa9PFukyB
Yq4SuLXPQ/jA464Ip1HXMoccDktvX6Em2wrqO9MwTSVTU+NJqxpI3klfCsXwy3Bi
dx2QSDdw7LBPU8mzvTUJXFl3Pia9AbuRkrSjNkOb9xKudjNbLelI1eayVbh/rdmL
2R3iPKu0MgvdApXEKP/4qY+b2BGbYXsKZMFg6tHLTXZR6zUKf89p2qqrM7pH+E1x
jgE/attc42qqCzLtWSfTBq3vmqlCU1Ah/Iypj/dQ5Y/BQS5vvP5YioQPBGhDVYi3
zIYOrPDXDwxaMaWN58xFxzGnNXmXpiN8mn4Y09OCIc5YY/gCgi9lby5svnzRMYZh
kzzjWHZpX8G1SEuBDPHu8nzdwBeICVV3qjNLDwvEc43IwrcZdecKhr+rWk9Xxb3X
yYNTCiD2OoGo6Eg5fR3+F3YB54mPJIlzsBvIFhGQMUv5vxiMwcd5Ydvz2aeyCQAW
rRcPHDLV8UHvKQI2kieruYWSHe/u7RJuFoYPwmCfSr/DIN05gdNOpivPSGF8AOT4
bG1jWesehHoz9ySPKXEUfb7e0Zgwmi8mlPqTqpdK3PfGlbDCVGVDCt8GS/H58cF/
tSAK52O6XJE+hp+H6qnIpa2i9Z3NJ15lxgD9oG0HdVoK6ZsJAeZXZjPUcYsHhVR5
NCE3blsDcZIJa/0wNdWV+HyO7FgwoYAS/iFN5C+UNlW0nYVT4wvdTKDRgjw7fJVe
DC0PvC2zo77aqZ74h6qLoxGwFHXIPuNElsJ8tzTUKdzQ1iE3N9F7OYBW3KzaVk7+
QLGXTlaDAjN13SnHsOV67QtqyDTa2sIXqrP1vOQReymylvMVfPqsyQ5a9cp5MToA
su31c6KrYEyIM8g2wqfMcf9hnv1N6JPixXy1xdj1gIiiS69u5mcccPfJdjs9RzOJ
B7U2YuPkx+LyxhNJgkTHzq5PXUP7oIfbd7xSEPBWS9MRzxg+Us9C1jggLumUuE+6
NAL4QTN/Ofkkh2Mzy8+6LhwHcQzA8hDMsK5y1bEHjK5ofTCpUukQSlwStcwRuSuq
zh2CnpVm/Fcyy/MutQh1+EbEaGmvCe3YfkARloAPEy0yerRYSZVRLcAyt+hQB/iY
3LsgORH5T8DzZGle7bf1G0frCoKl/GwtKLhzsBKI4mRApIHulxZFMocKbnrVv4q9
bPb82nuQstpfrgxC0SHYc6s1ionWI8DWzIv9lcWVN41pZS7LD+gJsc0vgoPDv23L
I5FYvq9sW9bfHVr3MepyFqTTjIbnmncbbt9eTpYI5J7GTCmZ1LZbUh9ok+9PPV3u
aJLRSunbe9AaPdPblgKYDp5GTiuEa53mZZ7Cj7xdmEB+rBwWmI9GSD6VNIwh33JM
0bBaqTi49vngpXdcXjumCnfVizwbWn2JLbSzPZekIFkH3offuVCaPasE0DtZbnnS
JFtmfLyIT7VumP0Oi+yX5Lgu/9X0kk1VDJPU2icwHufb5axNt2aPZc78JLFX66Cu
9fGpIb+NdxMzLWwalIoB7xPxF9/Yo79hKBiTJQcAc9105HGwkIHS9+j39v9Mxg02
MuOZHL37+Q7EjAwQWgQbZByh16GAYZzCXHxVw7mogos3R38wnCKbbGmy3KR+Fzzj
sSar+tfBwSkzIsxopz5WA3b0tuM8oqvGNP44/C9j+vCbhiO7t9mfx1bRx6UbznvQ
AY6c8fw/uS9yLr1gaQ1LGJSdOZgXf7wea2hOvvrifNfJp6d+KC5eCwk4P/+us3SU
/6SOB+KmGpJUj27T5imYKXp21ZIDBwGFLNeYQ8rk9hbnulUV4aNEL5lpKUG3pdGb
AP6xTz+XUrDbblBhqeI5WLv1lWfbhvDG58kdSgpHSHphXYNJTLcXnwpJoQgLz3xy
gIzhXriRqTw6iNV0vJJLumSaEAZ3iIZeM6+r5p/FYUifaXcaAiU4I9uQ03oKF89b
axvlw3dUv01Zrdabea+50g+EPTZdV17S8pY2L7CVSibJ9E+yAL+y0Bgbu/cVnZdW
Kwlkp3B0lIi/6fihM+7m6Nad2fXvcraHMKSvXEh6yKBDm8bwc7kivdBNOLJYAVr8
GO3/l5wNDuz7prnr2MT3AfH4XanEoVsnp26qWJ5bOpyfieUQ1oLPSErYVUG9C2Fo
H3x3r3oj+nBKICEaCrSW7RX8Cn7RvFCxF64FKVmAcVDRIb6jccEXGc7YYK2/QDhx
2Gc5txUKi+pRAmaSdcg+PR9VPPX6R/AMVUm3IggrePw+c1WDA8PaXv3HVqRfHzPB
6DCR13fa2FKArwYGBZP6NsrNph0vfAP8DE20gHpIOUbXkkPh9WIoJn1WZVH0XfB0
9l2zC+iSyezfIwjimNxeWqaOsNK/Mb2yOZf3oQP+jcjiasOrL8wzToc1CyAgNi5p
AXcdLMLFtilKnG5lCBwJJi1rw9r79yoaXaC4TkzRID0l5fT3f2/OSeqB6dMK3g2w
2en3pNVUVZWoK4ma1xXNLjt7X7+URQ2uzNTecuZRO3DiSbDvENUL9M4yDpP5X6DM
4o5/XUkfPkEYjjJEzeta6mJaeeZt8clhhpzMncugNVJnGyvk84jifFj2IJBOW6Fy
bIPWTmnOXy3anGpesChVaHtYf1DlOZWzHx2+49BtotT55ljOhkCwLOPhh+T8Mf4e
/+1pilyvTdsT1f8jo1Mlmor6WcxekyuelCL3q+/BprH8aujx5E/BA7xHsIClYTGo
ZCz5waoaLRmPd9IJMV21kw8A/dbCjjcYAqWQHk4WfI2siKiTsPI5gDyKIb1Ac04K
PEyqvkwYAcP6JdLPPAW7rdtlKhfZE7736wqBympVvsAkXdzDsDcuJmbWaoNZbC9W
lMK4ma1JW8/el9r3ZVEql0KKAOLI6HFUBcE9jvPX7z4r2cyVKHMUIc8KanL1H302
b2mannM+3sgz5sQ7iq9V+/LBrvTUPM0NdLckJ32UUY2mvFVSeLZ+65KCYzOxlj12
feQpEAeTFHJPF9jyfiWq7V8YehiEgKhuoFyLXxmmRVesPaPMQjbUpugt/QyOED2K
7CmqmNfsJbKuo+YkgKNdCE3eFxDcQ4ABFLwoZJdzJeBCgwIqs1UfkuekNSHeMfB1
vLkjFTyFzTYBvMq5+dTrLv0n/Z/kswrCYINXjC+vaPSH4sBB9Ghnyfs1XgECoQim
ZIt01T1UsknLRmDkG/yS4JTPhpcUK531+HfeOEtBvEAyuBZ7jyRSfmPodtkyBUub
tJE2HVZqBHNNdAxpfzJZUCFLliHj5ROi7+quzGC4mx99Ec8JOpJzwAjmjVG/yhgP
8QfEGpNbfHAqFzeYozz6jSlyxxp8cqHb3b1ldwS4j6c4a+RT53qHM4EvCIZ/UlXF
XOwqpYNptZincykpyCZu5lM77L3J+eFHjQMVV0LibrowXUjj+0Ep6fKFh5xS0icA
n/M/3sTD035xg1WIAcRC/Pl93PKc4rFQih3YV9kGxnDZP+nnhD2+b/8PY9RrT+dZ
HL3384FnUU89/mjI98qa+/mtquWM0FLm8e2Ztnxoc6Rzw8laLXMSYXc7y07RIfP1
Og/ojeySH1KKbCcTh64OMe1Xg6BIwSRSiMjofPd3b20ogAa1L6feReBURo/EyyqQ
eyBHW9ljbKSqh5gl9zWISmtbx0Hg1rG0L+yiMxECDMu0B8mJouhmtiC9lugQsUOk
QcKEw8MgwPIRyEDBsywCVVvd5viiPwXBDOslqqS+aYOKVz2aYmPLFQaYRMldrGp3
QQiIXIpSUKX6YEBjDrUe1w6FRhzuWK6qRy6MZbkuxvhtAmHWdFCJuyzvCgckK2o1
9pxCsSh6K9q72PNdOzvRelO9TlhhbC22a1UJy7AuDlAPbajzfXRvbPXyU84ckQ7n
XF/irFn9Rt+5XClGQkn1j4NrDUUEcqxK3dFiFMe0S5ERuLV7799rbTO/CqRpLaWA
1qf7zObu9qpgOYgEg2V8dE2Y4/18XGLOJC0lxnUD7uowd4BPa5AObLk6GQtJ6iXO
xJW6X68J7fRu4Gh4MFjOemxZfl9NNWyxRf3jVX9/+eWaXjUPfULvWFJRPbsPGaul
GUcLpJ3ABWZtny4qmzFboFw6scx9wIM8kGAhDY7QAh71mVYwVYX8knjk4nrk3ckU
htDxRPG+EZfaBxNKb6NLYyupctPgbU2NT0gMj5mPAGFDHp22ybVx6Cq1cCgJ2C70
42GazwvXqtHp+gow0taCJzBxlqH9CCHyak+VJAA01w1JHXOoSy3x7DQEW2G/nBuR
Cj2riIpLFSd0Wn8PyckLTf7FPgDhw6oj26nv+EP72Z7ce4YMG/qhaJKzFxBhofdn
6eRShNDkkQNDtrNBgVda++yfigFl/34eh/RU+u8fYHfz8LemSW+u8UaIfTAHt80S
IROquWONVev1sOcq18ETEv41Qko5B32lljHDw3v4/0dwepeSsmDPtOdwf7xEFQGK
e/eBb3Z3jnXIW1ecq4ayY8+C6coI57T6ebU/lFXGf4Y4SWS6833aXpu7qa5qAEZu
Vf0zC4e8602XozUN6uYFFCuDrIyaznHl/q175JF8R8L5QwHTZWN/TexnWNbvYlAI
S/050RD1m5WvOea6I6T2lyn2vE8GUFM1zQ3+P8wTsYyjzJmdiilpGs8IS3HIYLiL
nvaooyPYKLqBtrtS7GP30MKR8Rn7r58u98wO2z+zK12/+1HN0r//q9LJ/D/yKA7P
D/bgUpX2sCb+7hCkoumcjQRu9PSXu6XTUqftSaYptBqtefzXY6BmP4qdX8Rngk0J
pAUJazpgEziU0Jv+mDhXm8Q/z4k3lTd/1cjr/UTZ7eKrCbMscYkadXJURyAl2Rcp
OVYw2HumuqDz8Sz9VJgQZFpkmFJVKXJNW5rx5vtft9DbnTEVLm1cXD2jabKGju9v
382Orden0RFOxL/duZh+gljLwAdg9guS3TbunTUAJNaNNR4kc+Q2rm3JCTp/48BG
CR+p3NK9zWAt6MiueC3r/7RoCIgO4bDkgfuGWSwmvCmtPChdeRGsYWKlFHmzPnBT
BrE/eWRfLfCqq5hUPgYldy+JtnOAT0dr4P+W/FiP5x519xlaeVK/X3FDuZy1Vjb4
0Bgw04ktmz63ZXCUIa98DbFrZt2k6PRwY5B295tMrQDS02SJF4YUvISPRrrdMJK2
2E45zmgQijYQCqZSFtMwZlOPF+WneJdwCsvV2T5Xu5U/lBdvc8fheSawYs/B65HN
UoAWI9fIf+7vuru2s30eji/dHFsJKqPU9xr9zxJcYKbCCMumCLfvxseRpvSoXRWp
8tdmMCnqmQNX6tWRv57F0hAD8L9vwiAfi7+bmeOu/8eM+jCx6OOCxNfj+7FkEvuC
A6Ioy24Hx4xy58hf3KeRzC9nWZmHn/2OlsKNQXARCOpwpIiSgmiVK0QKowgfwvus
wMD1lWzuXIaOEtKonYQGPmSgHyf2eZJ8eI+P9XmqqiTX6Ovb7UgKft1Qtvb1VKDe
rBwVX3y6n7sU6T8Q/9YFaN/dgZpWGmJJvbKq+KslOwFCelz5vjbowVeDS/k4j6SJ
IwJildW71wQUh45Wahszlvw9dQNBIOZXFB9ry9ngB2wEwUYdRj2XQ7FrhZ4t72P1
Aemu9njlh729P/Y5p6fYYY+ubbxy7AzC4E52uXzeoqdcpWdaqc+PwikTDWIe3zeG
Ct1ZsCCF3mILC1bTLbGmCbLResxl3uQNEZB2iWRu05yNayNbysOzmCEETo6+BGav
GvKcgPIF89ub1cwpJ7LG8Mrarp3cDfqo+B3h6IE3jWvd9tACZUKzYlBZ5QXXUFcV
aWRmTwjb+ckttTsFRoI0Wve1A/cb8Ly2HYmNYoQBCfNiZqR1UuQR/3y1Ustk1Q88
/vkcYh/npfrgOZNrT0GrJ2oMCYkpv7YR8sd0mMgH/mUcaqWaI66O56KRNEKEWRz5
VCdSp3eQL2oFRIoCUcmh3Jg6cyt8L7I3aAObZQbHpuaSNKNF6hpbr2vEyVZQQKUl
9cZzP95GiEzX/MkaseUbCQ/T6P7lLEownjvVTugoMO+9hyxoQf0anF2YTSv0mHLY
by4g8SYM19NbJXIjhFeLxCi0lVl3x/vLPxLsXZMl2vy68Lz69qfviVxVA3bw7kg+
hCifmSjrwXYYJVzjzMkP8RHaTMKVTukkYvrPOkxWxwEAPgAC1hAeJndXkpnC4Dxk
hdI5E3krfUQdaWuAL8/g9mQTgpvu9MuK4IVmyYPSzkN7fhuUUKA0zkgh+sOm54nM
lm9BWIelhl1hL3Y9PmMlwBjFR7MU98FQWkw4yj38u4QBb8IA3mzxteywwoNVaXVp
R5Qrhs9v1lio5zWCwh/QvMjRzQXcN88aVXG9Sv9GSOq5/ujEUzlXJHBCPyiX/mWT
Mtc4zMAbSKOyLA0zQTrzVCtstBXU96U697u1bDl0rnLYH/GmTZAs5JOrILk77nIA
AelRnR6f13u5hKOIgXH36Gg72cxVLzrWUeTRiNOTHmd9QMAsjkVOPVGmg3BlIf2l
F2jj/68AFu2fVy0fgRE0BpEKUzQR2ft0UGsP/kbiSKzjhgQ3bOtP+psXx0Cgjyio
wBWkQHlWPHHQB59IVtRZGUYoWKbS/iVQa9xCSdGKnTThT76o8dCjVbcD1NAKTIkx
D22gZslqw+WR5yQhzzp9ax7WndhCqo6nbawVabizIhDU2mFT+Lc6zg0vze7WIRQx
tqeLZJ4BellcNfkh757JwclAG+Q9DvHu6zQww+Lb++3R5HL06Tkp868R4dlV+Ll1
QujaOF5DZY/WsM88AbCJn6AUcAp6qrck2JAikA3wwwNZYdwyN99ycU/tp5joL7WW
fGW0a9HioaKWx8BtDRiCTxOe5k+Uk+2OPQYmOzHjaaszUgCKDloCDZYKpjqiMGYm
7KGMrZDn2WktHBQMqF7VCmoKAp3y4wEfX/n0jUnf7M74zeRsg2fBoCiK5sVwm/1Q
F2+wbES2VsXvhVLNODycdVpxxgKN1HEUAdvrtYgVZbqLySUPkODCNcZVcOQ7lu94
wEab1S5e1hEqUe6aw0BWT4A53l9g9wzYXuTMYY2bccGAR/3pZEBbLJ4nul7bYjcI
ZsV1jOhXs+/i89yb+Fp78LAxSvR1mnIi5nSEcfVXO9sSmmrvTS7SvPY2mFCBfAmd
Rwiw0niNsyVLQyLRxCGRhNlT1O9QwW+z8ty1GL65IWYM+nYvg48vkmsXFqOBTl3y
MjTrReGF0v0TqBdJMiLtEb4vQKBMbVSW+gjT30iQVX4v+PL5Jursfez/t+4flz9H
gH38EGVOctOB0B96NaWGxz1BLN22qfj7qT0E67hbOzGioZB6i4w6rZZU5XQ1y49G
l0T1dIAax4EYfdZ49DottrFB+MbX4mRk9pIpTZifr557cDaoox10ePB2JMFsWqYN
WIX9Tg8MfotLT/oLhtMD0z4mAz4yaVGmRUF4VvDmuoTLcBXLeMagYDVOxOzg22ia
JywayzEqbcEubjLxtrmRgEhaNaZXmM0jFGWWkIKC4/SdUhAplANQR/LxDFjVtWRl
DTr9j0U/8dnaiQTWQivYO/NCRNKjSI/vKjT9Ni0HHpVM4007dOljjvoCcpBsbtU/
BkAEmo+CztnepH1C/IHt1RtbBv4j2wpiDq3OBn6+d/ORC5v/2rjWBQpQsYUKCuR8
F6uytRdxgqEJGZ28VX+59jE9KhQE6GMtC5OTeUU+aWizyklLeTSmidVaOqHv56GD
pNcw6uN4fSHsrRITTPKWDcpzJm6UKJ20Gh+JOYY+kcuprVQKsvVXDRlDxQh34fsv
Rj/pm9k8KWMvTPh+EEnyMVNRtxhnB7W0ow2VtXBfGInGerm5xVzb8QjOEwjOlG9f
elTdMisfwNUTdGozcYb3CR4X4SRYOwRCIzObT9byzGBA1RH5TSC/S7ddLQekxdNz
z1OSGRshz25/wRdCuaXG68gDD7oP0ykrOrhENQRqxI2Lc1yBdzgn4SuAgPLhvF88
j3lj/ZLTSen8k02BsuZiBqnZ3XUO4h7mn8q6izKZeHB9hiUCnpFBg1/WxR98DMh3
IwFsB0/c59O7cxMIcrCbECUtaxeqcvDBD7+HQxL39XtJb6LXnTy4WAwH4BiulySy
Oo4ReXyzbVY+bIXEFxxU9Z5AtGH/THHvEe/1qagLqeGcNp+jYnrF6SXEITcvglfF
2YWeLEPj8gjZCBSbiUEK+zaDYA20zLTDzMl/klEUIoIOujldY8QhtBUDVS1kvXej
VPbqygAlfVR8m3YsTMkfjg6Gd47bPZLr9WK8ozl1CdxoE2GGCECKa1mziy4HpKXh
uJR/8w3RzXCVQNfQdwIGiiYyNs8ZVuDfBClZaEBUKGdfuPeCKLJe8No8jjhRsTHP
xTioLM6rp60zaoCBNFg0ogXdGB3foD4inwgUG7yXiE7BY+MOeEqIDRFqGC4cW/5b
RItLbq8imb3Bwhr4q5fZ9kJZKVuzOUd3LyypwuR6r0HKgaM0tr8wNO3i92/URXcO
3lk0A3qYYBUhJpI84PcyoKFcBZ85zzJBgwHksNpWvdzBEFtrkK3AaP8XMqp7XBoj
xVSKTTFazshQ1+XZedVT67pRY7U3yvMlyYcSdY5QHr8Ukbl6+5LFVhKVBkd9mlN+
ftiOJmPfqGsgQAEqVI2v0ZirCL2YOrEfBOVZO20mwfBR2tRwF8OIaAIEoOC0hoXT
V0btztdppkhVkVu2RA4ZrTJJ6lBGSdM0ZRjz1qIZzLb3do0mRflAJto1Wo5gKeYP
1Z9YI7HB8mI7y4+5tOUKBx2W1JoKJQpdWiuQgrHwc45YVTI7PYZWevCVjcbkHNp2
R79zcYT93yL/YNagAa+/kKjyllXk73o3jVjZpMbU/YLnP8gEO4NFCgx7+HHunfj+
1pkXL75vT6sA0W4GdzCTU0B8Pox+sNjYNSYXFcgIFxI91Zh+jWu9V4x6mTaweMyN
WW6ooZTKvEdMu7/XK8R7rMSqHQFO7J5dKM/Un2vqvMAW7MLnaE5opI8hQEQFvYA5
L4VF1j/HA22OFrr1OqkZx+mGZKCKahzKb7xYa8cXgSF57KU2mJLDpYm+j49XdA4O
3XgYCgJsWpmVh02mnV53hZpp3VrBAa4lGogFX9iYdj39LR2lOsyAGJtE1Z9IA7+9
WmSukyXDAr/rT+FgLQ5tW987JUHDTvRUNbRAJ/uuOA3d8OfE8AxO6ss9RSGjsTsG
m/X5otwLHyDeR65XgWvpwANNsUmKjwqzgDBAOgbz4mE54L9Y0ixMqNyzjmtIyh/g
E+wkgv0JFpLOLM5XFxzL8wIWbHh/HDq+jwSKYjY7Jz1P4hLxqnqg+B8bdDxAqgvA
YUBOvI+TZa/gJAjxiIRWUqyzCyFkVThpl3ZTkvB50E7HSL6t1hPi9la8ZkXnaz63
7sRuQqo3vud875gC8yS39d39j4HQj+MOO7X/gNiXwrRgI9e2yUYHbwEIAX4lElzT
d4G3ZefWtiNSUkXCn3S1KcwF0BtecwR7D/GoSV81XbNhPcDoQXIxwNv75YnYbq7H
DkN4Tcl+W/+ygBZIRki86YHSvmJ/VEm7sHkoSwOhaCyAwWkvPPaGS5/CPhXCL00x
hHqfd20oJwKUHKGhyrh+1kqIcxsbLgFAOo6P7jWj5/aMlFwaobuXPCsNa8KY/a83
8KaoPndr4SV6+BHT7HpPkoLthQPNWNpOxXp5M3Yd/aL6lMeIG7Pf6gYbty82jboW
EZTYBbwiH0EFJhkprieRbHaEtJIZmMZQ3lQ4SRMy+sdaUvxeG9rxD30el/JkVUNH
5xOql4ZrBQPJQTp/gX0147t3GPItDzg2u1Vd07KSbl+7exs8W4KSoxNeLwFCAdtp
GKT5F6tiQK1S/nqKLx16GKSjO8hwZqKOq1pHd8dTIravibwoNjjcKlYKhWqIqn+p
o/YhuW7SpXy5Ui+Gwgr8KL/rkAcovOv9tgJJu70Y5dG56ZM0o2HJ3XWsmzBxGWTC
ZItw8JPCFKpZiddXulFTSDNg+uGg3w3vspIAwyNX1DYhc6nq5Qp2hyCa4P+DB75r
daugGs3HEs5hM5p9jpY4MivO82B1/07qw9uiLRi/tX6kqieExz6npgaerE6dCh55
HTwlO2qO7tcUyhKwkheDw+84smiY4lGIKq8jOf2NJfNA16e5kQ8faIUUKC8W9Twd
NQagoK4CRoRBtNxqwPGUTNntcjr76byk2mQFSJeJwLPDx9U7KbHNY375ECQJrY94
RYXjTu1SnqJBBvm5xISo7ag/oluFhKeyNw4xmYjfOS5oc4G5ZXQWYdw6vvKbv1HU
wCxuH22Pi79BjYgrXHL2Pfxf+PUjIoNZ9VaOPyY3pZPXDR+zky9lpORQ/TPTQ8aR
d/4w1yPBJr/69vlRjGAQo2TCcOdyQcIC7LIvboiTEEo9ovRlff5dv/8oTpfxEay4
xff3Hnr3AWTTBDuv9VF1bYQ5syy0TuKSOZlCS1sM3/WE3DJekf4sew0Y3wI7xHK7
ve29Z8n5SnodBhTejs2GdVs4/FG2q46EPI8UzK1E5wnbOc9RNyKi0BnSIjrv+aAV
Ok9Mc/MA+8fwU6tnryOcyuGYL/HrW4XAtr2/GfOSUSt/nAgWRLhQIsFmgmOcUw6Y
A7TtQBZ/N/Msqo8xzGvyhfouNZ4KbEuggDmTKMII0jaA+ZHwF3TJ1s6tK0wTdoJz
StcDOlc82RgBEWUp98QBzCCv707qRRoyPAvNMUTMSnLslweOq5E4f/uyvtzcAobt
zTxAwtSmwnpS0HZ+yHrhy1p8pW9pDXfoaLq6nzukaP6ZbdSbpkz2VDHefxgMIEiY
EmjOBlurzQXHh57f7cEh3gGIMMcS1oCp+4GwJJu3iY6nxTqCAXr64Qy4ExmfbvmQ
ZsHiBX8jlkxgdUfKKPSyRzhhPSsbNjzc/cNkHGpdxHmm0sU18+GhRZKQ5q+8AucO
9YydS0YyAKY7+ISgEh03sul1mfh374wyxdBgDdwqDrRUiCvsHc36N1pDqQg1J0hg
MaYm90U8TBnwVkZ1BGzAfSEp7saZpxz2ZuvQUq5KFHFRGNa1+Feoqx6kFWXobzWb
uyOETwKL6JCzXd10OPxGDOOfjDUIoTM8ZyuZ+hbptmww1EbpejiHfuswUcRSeRup
qnm9GY5Pc/ey61x0o7m68Zcr4b2q9bJIxt9Cno21MVivdlf2WzGIVtizWWA4MQpL
dpdMfP07SSF6QkQhkK2PhoEbzL67X02p4DBLxQVcZ5Eo1PA3R5SIbh2Z53u8LdUe
H2E7fTxt9OhYv7inlm//UdMkMdp4qOmQMoBA6DfeBN+1S9LtMa0UPpnrsOV731ye
EraVyTRGquIT6a4jefd5a2nNOnuzccwkmBY1XUZ/lg7/GNHp81cDPOzZo2a46BMj
Db1EyxePKFwI7YLezyxwwl9jgB818TSx9WE7qd2UCtfK77HIkSuJrkIWwD78UzH+
sL4A5u3CCqm/gTwzHYQXQAP5UlvFYPcYN3yfgFn8wSuZ/CFG3PoZ/r8sjsUJEMpn
WL35MQYAVu2Fi5cJJOQBu3MpoRNAxx/Hp7msceOIuhNTPiRzMssx5m2Y+NYuQq7Q
4offWCRU0HFwVmBKVOifuSAQNH2hf3K3emnE7M4r/WrhT6jifseq5Ol10WsZfHym
ZKXia2bAQr93skscz6MKb1UPi/wllVuVUfGhzNwakvKPF5WMgZvCIfQTVxYS+6fh
EBw8ttzXtspClLtePE+7vKXtFMqmY4N8JpM2djcn26Z5rl3/iwVVVmHzSnKFlFmK
TkKK/Tnrf9lLXreH0+hDr5jpSpD2SmrPuJhG92lGyiwBYF3OYCpcDtdfQDoUlyar
q9JyGXTRGsVvv09pSLXYJTYXSGagVQSuli/CMfWlYc508hQT3JCpJG9l6lt85RJ+
c8lSafF+FzFDkcBLrEQbLrA/8S9WuOmGoJ+JHOSUzs7IlF/DcLmzaHyw6bTI4BWe
NuBAtO2v8S/GiM+jPcwD0OG75UJdIFJ5BlfVp8HyI/qObUZ6tCkC4ktlIYmpGztz
HPETA3TWXbllD0k1E7uiyaKvl8XgoIDo0KRrBvE1orHNrD/wBTz0gfB+KiVcC7iX
RR8CnfALbF8DH5GnNHmDn9m5RpTclX+OSOkVG4twfcQj0JT6Haja7BDNHkk9GV7J
LU0+QZBcE58rYIkYPav/90qBiLInx5Ipla4B9FWgiSZ/FM+73kWWrPlXPNAw2omP
2koxLJ+vXxM8lS+4JsZoXJrXlKwwC50AdnPM8YTYGA3GEPCQ2oFBrpFGq/6E/8So
k19kP/vY0ukmTtiKA21xrioRLa4OXZhAL2SXjWIdUw8q1evrMaJGjpXzCiN6AcTj
2ErlTtU4KvYxwyQaPGXLZRJktlJ/PjJI10R3uKPWMwRA0T2Q7SFnsl+BRlwMc0Rl
qoeU4NMYNz8ted+/wFryhBqsBdFo1o+EhXG25glvBtZHxH+0YHphGB0xfquYA5DY
78/H6kQ6yE3Xsu6p7HdRjKSNCVL5gGlAZG6MV2qH7OMdmNsFS4yPHYGJwhVq2iqL
DDvcy+9DgiHNeknJKy7PkXoV9BWNuLWmSJXt80PX7KGfgfDDiVN/6GiBdxdiUYp9
DhWIT3N/qOasxtvCO3sIGHUyeH7/mBI7jX9vMRnGqwfBSZ/B2iPjNCJDXf6Dy8+I
ljew32CMVaH3xIuJ/+v/JbWU7Ge/UTtc2lz/D2KwPkz/fEzkNOMQ9j+LMw/eIZqC
VRiA4QCerFgXMuAkPSfo8UCNcnvgkBf1TANBM37fpdfq1RzyAiWANOWe73lysMx/
cemQxAdoa2TiaPxC6ZJjToz/b/609arK2RHyCRQWvFdUI9HgubnqEvPN34UXZnRq
saEvCZu3w8EpcAlzLFIaC/DADHhactwr3RkEUGmtlhs3oEoaq5xtOYsTpbtPU8y2
KhH6jEHcTAJliCTN6lDzDOlwBzLtKNOiN6i0+kcOWRjG1jzW5NxCzuTS3BO5C2tn
ko4uUlURzBWaszO9qM9kmIt+beCZBUVtQV3yrdBeODxkIvX/euEbA5JKmO7GQeNS
194liqmhjSQgj2tQSJWG9wfYoSvVbfIHGOJ7wvCV9YYTBnbIkCAK640Qu3sIrWQG
1Rx5/hxhpgX1FnTKKuRudnNtlGeL5IjNCWHdxiWERylvqVF92O9YBlpleF3zcj63
l9i+bIim3hk05p7gziFL4lrgYd91XQlZQRZpOh+EnQiW7efNdUOCoLHghlvMea02
2HduZPYj0Vo5XK5jQPE1d+zoMkIkQZ43N+fub982Jyj256V6EeGSYpSMxCvpZ8No
2+GWSksVIEU5PnmXOoQGpXnnWJXegH51HYIMPVThH/S3NPmrknl2tupdyqPwd70x
VkyP6LzlDkt3wnZteLCKe13gdSs1kg7XjL2Ob97YXxl/nF1eoiTwIAfOm9o/+OMJ
3GThYQmBx63y46O5AHloKor6kiJCQw+uEvoajzBpawF+v8VS2O7Qts6OjGPBU6wD
GUrMgYUNL6U5QoMk/OzP/1QAVbRN8GkNGtTwOHCvz8aZ4VSMb0wMD//IMObC/BDE
s4+nB1VhzgVV8yMwP8vGAA8f0ZdITBRus6kS7iRdHpPziHGiAjEgXvmGPTCMJvWd
szyr443o1XkN//RCItpjkFKPn3gmj9etyqS0QtqN7KDaYhi5MugBpp4dGKWh7+qw
cOWj3f/zF52TlZ2tDxfcM931LOfWpDuoPmn+lgiErHOOOi3PJdWsu05DU6nyUEMO
YS/zWJNgqDII4xOGwMn6Jq5UbstfZsBaDH1GMIy7x60YjT1XGr9dlk0yR+IYoXYy
5Iku3OX8Xz072uyQGnzGQ1Dpe7IYoSFpmIDWHeRux5lCGYN83GXOhDffVSjudtz7
TKbLZ/kHqNfxVeYxsvvPb4mLFbj55qBsTeBqj1JCmpCldfhhKl4T/6CLMccd2xoh
UjUVn3b7A0goushHuCitk5nt746/GHqXHaKy9KldQi0ppyHHawHKo5nZsRQUN9Qb
yNBGJYidj39iYZs4zi4lIp1bxow5PS6e6OkzGZakJ5sfhsYf0JQFxWlStZZlTM+Z
JbTGm5eeT6ueBqTqyQWzWP1hrbA7FUQVHD+Dq87IpCkWYsYn+monk76wDVTg4yd9
xflFr+SbnbOWXFDe8/HlbMTEniohn7M6MacaLfqc26mvqjqxx3WMD3wyLqEmqt0k
yqyW5Fp4FLNzwrmNJhDEPKByO3QPuWeoNOYPuEdmH+Ji4ClvU+nOZtZkzem3gp/D
Ryl+3xlvM5eHLzP/6qLDk15VlJm+Ff/LP9UMygh2vRhPU3K9020iV7bEXGZkNjCk
7sdotvnoPzsxyNMrgORJKhgV8PBoxXr3d6d+HwHp+AWg2jtalCZ7SepSo6ZY3M7g
hNPUqHB3D+J9kGgtZRhUctOxATAaZPl4ViLVIKXRgs2hRDwZn41q5l9dirvun5lv
CI5M5JwCrb72Z6gXFzh1aCFP/uxvifVqBJ3lARMstU0aMZflb5Rf8azrjXnNyV8I
GwI4IaMKJexJW691Ey+0goMKUXr+tt3IVFcgK1IY8mmKfp6EjMvy1S1zVvLWDJW+
lb9Fz5dSWRblLXDXFl7/tC08eQ+n8DwavLHXVBTe//1dh6jdgpbNhJwd64x3TH9C
fne17+lz90R0+UYI0ZSSD2XtahocnOs11gqm6LfJpBF9NTDgyR/eAR/bFv5HiXWK
8rTOgyk9zk782g4+I2v7oJteamCP86+B/HYlD8xISXcCVMKLgQjo02X7SBkWNUCO
YsHg9iqN1s9IhYItq8ww58NYlg36AvIaGiad7pfrKgNnY33pGeQCm9TXrm+MnJOm
zsnohyShxKm6wwxpfpSdM9AFRzsfnj1p+Y0D2TRTsGKkFHUjKPIR5PDI0BdtGq+A
1sTeIvU1WKxzx0LA6lJJ9wWOCO27Rv8feStkKQmBQaWYLqRJqVyxKpmsmFKPOUJO
c3R+2j1W2NjngNfPoHdN4FsfCZrXipgaOj8N0wm4hcErj0uBhEDJ7NJEAKJkmxim
WmIuDvKnl0olmgPe3JKud5EOUohH2aAjL46Ejmsj72IBq7vNRnlmu8dz1HiSwpG7
8oIh7gjRhWt6o+401AxKEhbvhkI2Lvauwglf38//5607YDvgVma7+dXlE0YTTJhv
eGA5ZbBZRvzv8ecAW7y+sYpu+ZojzRhqG1Uj1BiyPXdN9JsfnWG9M/DQUBGXFn6o
uCGlYTnC9RwlSshDxVcORk0PMdGHv04NuuBda8C2W5s/qH/QtX0JQylp7a86P1P3
cUzI0YU+1ki0JwCHkWCqCerr3H8RnGgJD3bc+8x6qwxs9EfewgGo18+O9TYvdKSx
K8YnjjtZcUDxTP+x4UboUa7P3W+2EHAI129bPhIphCi+z+3ubv67dsUkRhFS87T6
uMTvhCm4Eez1Wo+snO3XtMA7JsISGk4oIAWB1pHuVidltPBBPmR4opLTsv0W/UOg
MxjieV6XdEEQyKpf4QVCnkL6+y3wbKAimrOZytVXaBHEJr2asMK1S6b0vJcMTNr2
df5rpOlzxO6x1pQDgbxWdw+mJeUZIoiuRLoKUnhGW7ej6yWeCre6ww8XfaLOLrgX
hjxpJkJciYiSnmL5iZImp0Eq8IH1c8CPAHVTXAXhuzQN+lrCsaJXYycySaYqT3ch
nGw5CT+/uz/Luml/mlQ8QVp5jjleme8Dq650hgKqFtsmsTQhSAFbHafxta1CJreQ
jmf0GFF3KTyCl6IpvGMeSsE9KOZejmd1NArUm+ISCP/2Wriq3y3W1Z/TsXEEFPFO
WBF3iK2c2WOZkHOOS4gNC89jpNrLNHQ259JOa29T/1zuFnGNL1++EeMqumPgtPfB
zcOl1zkvoPyXYe/EFcFbl2LQOSozzEqzsJfXPmmjXke/AbtF+UKwsxar+pPeeyhO
oq2wBo3afrOt7mlj47ZdR6M0qKCKszx0dXBxKRoCQGQE43UfyS8lxnHcoeAqULUB
o6BO+EKecwJR/AzmCxFZ+Okc1DYpaWEKHavfZ+bv+zo4NoOjJ5Za7+qEkCOxggok
xTYjnu8sQji2wN/Gm7wgvRG+cy2ZEldK8eesGsG5HJhVZzPQj++VhlI1xfxP9NyP
S2FLeaY6EpROSoZKhUO9Yoq6xq1ioeoNKkmrBOVejHbRxWNBrtIOVIhOhc0uBH31
or/gKJQQe+bJ2YF7kjMLk+DXksvPSJWIVWICtBrTcoiWBlczY2CGHj8YNPcIyJob
iOdN60vPO91HAxmyj790grO6Ql1ScR1ICCRPiCSgX8qhQ8TT2MZkFAESRKsSR7rK
EM21AhD70/bATamOhQa/OEbhajYtdz1Wd1J6EqmsZtpuSL6pwvHsPQTloz/NkPP7
M+XeFxRcUzo9Y9SDOQKm0ziOyWHkGwsFYHVw/nvbCcG3t1O+vpMU3J3ZbIVoSh/i
OL40MGOc2vhzkYCpZ6nWA4rhvOgfY4S1WSFpeRjULGAVNoqGuZSFtlaQSAEM3rNK
K6d8JYDeYBn6eshEfayenSl/5VxZ6pagmYqjIu0JOsP6qJuR43yhLwjFnUaPD5QF
CROilf45A/yJ5Fs3bAbfM0w7MOcChAScJ5DgrwbkHYNGX2UvUT137VY+rn3hhN5K
JEhx1/i0VxwtyoRaLNuDkhBq7q/7DvD7OG60N2e6txfLuWyX5+DXznrVAdNflsn9
WF1koB51WTxn85zd72Hy/w2bzrza7gstHRpbKp1OgaiqiDxg5QlfuUW2ntbjmG2K
mKNaVr5Bf/uYNORkoIFcCdpLT0hda7igoNp1/pF5OctzOeuOz401nELHkg/AUYg4
OI/XqH/PQBvMr+MqQ/tvpeKmtkHAumvGN4/aR1TVcoASKABQIAhWAhxMucu9x/82
j3avkM8JKTZfQ8JgLP0QfeG5Gj7BFAPlvjO5pm2EFnezamzncKoWZ73OfjB9ykmY
x8cA01ctMy89O/BslWQkSdZn85p500BTUoHL9O1uqBdS/mP/NLslAn51u4EzJnkg
bW4imS9xHXmRiyuvgpX77YiLwDjGvQFEvqhxkv1HFIrB3qOwkLXgd3LWNMZiSv+X
GLhIip8JRFBcvGawVvE/Bq3WtPQWHRaoicUbLKVlFBV2FGea8ZI5MMkh+bgGdXzk
sWMOIYsnb4lxZS7+yMWu4TtN01vCAv8s8J8LhiWEcmeaph+3w8Ls0OF0w52Yxkio
nJ0+E6MnAmzHVWiXBpPcjAWHWEpE2S5J3B+o7CVfs2UBvazhrRVqhkAr7wIkejYQ
fTDpiO2RUxv3vpOkurAw2ltibN7i1iuPsHixLyi3mehoNX1tMnEKkBgW20+ZeZuM
fRs55zHoqzig7AVJPFzP0mw2zcqatDeAHtvE9w7Rr3MwOMxfYxBtD5F49Ec9LDmT
ucEPcdfnXoks/5QERq+JdgYmAh+PZbRoG8aGklnpAyB6M0OyOs902bJege+kScZp
g39PJmOET8V6qOqF3t+TTY0BSgNPFJfkEBBIrGpp+haV2dIgf/gSNLB2g0mIxa8U
KsqZB+4FzfbS/Bw8dP6EfUN3HNY4OOlJA+1UT75IecMJlTu9B8OJIJpl1fReBQrW
9Y4tOi6MI6a0NrsZmRHm1kChSX5YGBVXZx3x2YGgfM3s1++yCAcrTiwlOZBkvex6
QhrXet7ps5HBtWYaOgsEA/BBckaOKCQYZQNYy3jU7tE5EoBnT2Pmpz/stskx3LxO
O57dUypvTx0rqwUMGgBSSr6iTBRNkFwq3RLSTQ1nCSvCrQ2w+ndGlHcL2da6p4bN
R0oifWJpuKp/fuCP+9ErQ1Nkmhh6ln2YEcZcJPKDN291RZSwguQZ8lCQJWestpc0
srKypBAyZ+6z7Zq0T0jWN734JB/KCeDQsCKhgHZ2uQJFImtKsG6/YN6QGOrcgiqp
iwuh/aclZTp28mTdM3mH0yvsyLpBPQtV3vddOTP8QNW4jBExlU0ggBQKg39r0GBC
JcAUg+EM00tFlJXMsDMAbmaurWgkAzo9nKmjfQAqaAzkt0eUpbsUcHv/adUUREGG
8q/AP+pLdrpVkp9K9HRh6HmL95+rVyobaTaTPFxmhPgXA+dwWC7iKhoM7hpIPLF7
5HuSwkp6uDPwLWp53zyFMj65rrucOXbprOX5k/TXlA2AvFMgFX3Bk9K9ZWdVdGli
V9Dt+i6jPnXeMCSDHV3lW6rbu/tfwAMPMGiUKhnAtSgkdRj1D7eVHnWSvNbAB5xN
nAzvx2rE3iInqTVsPDBJMGb9MHwFjVKEpvMxRqyF1DcM/HjLlxfC7hysu6UI1DOx
8LmfNRNb4t2BqSdg+vfeg9xZm/0WVREWl9A54l5JYRdEWScn82jRLA1R39xNiPMJ
6yzJZQJVnh/Ab6FaG/SJx35OHrkHUts7v7ArjmToUat6mdU5ZahhAvFUfFs93ble
veC0A+DReCj52Gizb2suiufqSwAh58iVlC+7Kf+p+0BrHuP1mdsAwS+fCXz1w0cw
lj60YtCsYiNEFfNph8Rmr8pGekpvI8VBIpP9FcJpT9esuhvMBW30NYpUHkW+gxNv
D1T1UcYG+mTVqcQ73S2y1EsNjmmtgk2q8jrub0KzvSfkQ87qK2lmVBS7YNpy02Dz
gNAjK58vIWOqzNRxlirR5/KxWsO6PtQye2JR7AhJVIVNBRR7EKx31KR0iiuFvqiJ
kWuE/lTxutb0zpyhjooL8j7GG2Fyuu1cYSwzZv8MZOEo/GjVHw0qIHaMGhb7X+HF
QtQwDueUQ5EAqVMmZs8RpsQpSQYB9RE+B4RzcjxX5YrRz3nT8ZxpH6FN32dicrsA
4oKvaN2OxydkOqiSvB/dlugYNeCKRGXkqH5Y/eV9IUVZYzhZ59kC3qSNtSjEbqH0
DsvYfLuRzLiRQeaAOl1Cqp0xg7oWE7RLYsYYlJIRQ96T2Tj5VWzrdjfyrhOThCDP
UnKgvqz6jGpp1XkYYIsCAJ5L9UC17DmWcuUVNK3C7jD1AL8aHFXNNejG+yUzkbmg
c27R34SnWcUpbNyKkeqZAyV+RH+FG5APOcOp4R8nRldDhdhgRpEv9AJ427zfaPuX
TZ5GcvD9mADS5SgqqPQWZQr8aUhMAs5Q0L3jr48MPdTlQWAsuEWbFE2sLZ1ZIQOB
KfhukyrlYHNvWlfivWIi+5SLzWVnoaR0zDck9pq6ox54OTd48XLkdZKVoYkBVtbl
TR7qMbSz1kKQVG5cjEK57qPmqPELwzQeV5ffQHPoLW9g8UJ6H/JOC8fOjU2OzuWr
WTJc/GdLX0fEUPkvqeVcTk2pmplDjV9K1U22+6mRV/dkDXjyrzBRxsi14hu+irBa
wNX05vwMj69Ty8ME6GUsj/mLSYAPK/6NZQsDXvDfck1BeCRXZcH8H/73LPSqgbco
XmgAuUIOI4nemI7EGGPopoq/FvmuyXYTkWWUnLI4QW1VAGxHUUEQDFBYHo52GbaZ
8Ve7zD32q8xmC9ryuctApseDoBjtAVlNXWgWXelEMTj5hku4VFVpBFiLWhs8cYfb
63wNsuEM8qfDkMibzTwJARgUpmgVtr/Qs5HWWqarf2VP3HtUbZ4nfkHx7LzyYFWX
RNbVpuvSyuvI8RhJYKMPMxbaiAwjwANtBPxDza9TfcNC/h4YdMfcpQHnCcezSaRq
we4rBlJOLkVh3q3IUavMiskRaRpGthYGn2VgSUiiCSfjOmzLoBu9AOkf5QrpD3NQ
n6uIqCaHyNtc1FgBqBbvWYDcNrLiTb8+lYbMFxUMW4YDoFvrI8/qDA9C1wbAXdwh
9iyTGbQyDR5vTKyoCbFFRK9v4SvG2Vq86CHwtmGuIlEasU9TY7oUiQKgrAUYV2UC
V8OgxeLoIrJeeuVL9poASJUP+lz6Uu0+i/1Jnh006tN5kZoeIQ1xsTtPI3Bu4XjK
+IwsxAaOi4f5xmJ4SIuTIQyIkvM7JeFAorOa5FJ2fFsaHdD4QD7+Q3FvpL/GndLh
x8O+eqNTU6n7lPtGX/KRwt+jU04P5R+XcpPqHGPNAUjeiEUavXlTB30taE/9biX6
ndB6b03oHDCjACBslcQX+L1ZQ1zBsZxEVFuZ1LoVS7wlgaqy/O8QxYAAlLDqZbiD
j8BnSMpqT490Mz4PX9kgpSV75rRcuNEH6NydqGf7MGQ4cB31nnNvepXCD6855OSw
szEb7i7Mx/BfTGWpDRa0tB0qdG79ZHnfQMK8lVlsDAeqAhzOvq+ANSGZasayuBgU
fTOeYQgkzQ0G51PyXZlDlO+JYBkjDbZsTRIZPvfzit5ewZ5SFavLwc07Vm2gawH7
SisA7xClWf7YGcjDICx0Jq05SzlcvmaA5dM1oiS27Ux0w9RutVLwix1JRA0vGPNY
MpJxg9DFQd3vjj3fO601CDkD9Wa1Ji2WjGggZA4obfbbcpUI3VobC5PkxhIG4IvO
sIVuDtkLeimgkeft5CnahL2FqQ0+9q94BDLIQLYBwTNNkU7iu2Aond0O96W5PYue
sPZPhcdqJmIDFOE1vO6c1IAChh3KqkarlAzlLFsaVkdyDCLB3CZyKuK1XGLH8SUf
3zc3CHEtImDC89yFAuYFT66EV+/wFi1GuxJJC8qd+o7xMh+4NPJbGEx+rr75Pxm3
aefHDPIO/MY+XrLfnzH32WaDxssb/UBa3fFLx8TsNl2YuHMWueTo47V9uK9M0kdl
hyfJzvrZIpUHv3a0qB/xj/pc/wfs330AITxFL7v0DLX9n0eJy/j2T9G8k/dlJEeP
KaJdn/ceQ+LWqH8OAu0TDwf3RJeiJjQovdHH8/rNnXSp6YQYC6LcdpjYsq+f7+bI
1RX6vsulp1Plm/xva/5HCIe46oj6l8lao/SCYN98YiiqppHGCsStR0yxcn8VXHeA
aOB96+Q56colOM6GcEq3vbe0SvLHDqwVqMlqcSQpym0lPJMWVKU1WL7WD3wRnyz0
YbSkKAa41zFealxvvuJMWXV4LKVabo/AgSrfgbGzx5KGYiKAG9vzgSfZQGNG0BOa
4r8EuhnT86WvLPYCkrZ7DfnY21oYjIYrcfIwgAhgLpPmEOGlofs+Y/ddYEmDx5wx
6iv8pOBAYjiYLY5hZ9s6E4uDGUJBjTQF1xr0sEWSGp7hPv+7LwGQgsal8gAWTIH3
gXph2+63bp2E1XiKZOY0bdmfVy5E/OSoFVvYkAbNxkQmfnl5DfhTiiiprA0rpZJ/
tQBq6FoyOdnghUxejfzv1Inu7kNlYOnqqBrQsd+6uDgv6iyQ55nAII9BLfRCO6bA
UWjFlrD6xvrNwBBN2Z5x3/DogPzkBET97TglVoZ9OdqQdx+3MNxjAxE6hwaXgovB
abNtcpyUUOT76W6NNf+EN1CIIOhRIdtWKclLzz0SINzpo1nzxcyWhq8G3Q9eHW0O
7jRcz0avo61ba8ybizaFOEhXazcLUFNB7A246BHwWsqB7aEdqhTrgBNJCqpYwheS
JQSoed61WG37NF/xjNElK4rNjRa55lphGZVNliBBanwoRlk4+kqjdzRMvopg23bd
7QysT+TddFiyCNtBIUqw1COiY1WFtjIbvbq0HMjWbEAk2CtGhoKCE8mokO32ddE+
lYUrKEfC/9ksTQcUa8gV3eE8rDIN1zoHZF5nPx2OHZG3tN+lY5M+gVjGIrmk36F4
eB/NgSQyoxVd46hSoe+a+pM2dSCXGXOChVjhZ09Gl5EPOOC6S7yWXWMMxgLxLv29
YkMW/aUKC8ZiFl9gGQGJSRCgJLYUr+BtQ6XkfKDAB8OEHt3kasPbo3O+E5ftXi35
8ir/5dmAsRgBOi+iq8TLn7qRoYZTclE1oT7+DP7kvwfDN580wC+hgt+rvUfwC2va
CupHReI58mglDSblIbLMCvnhQ7ROyhdKKYvoxU66FSDNjAowXhC3rDfwNJcnIW96
zfpwe31cowaN7qsQDKmsRJGH6pVwVsZS3WwSgyb1BUdlimCByB3yvBFNnfslsx7X
uCSiQnzrOKnkQaUvCqXkAhlK4ONYAYwZTrOxYnMB4IFsKVUjsvX3I7oRKdxSa6vy
cdQYkWlEA/KwzAA9Bjxohf/j+JaHtO4m4G1b8cgU4VNPzuEpAuqkwgpnBC5n0bCA
cBbi+DUurNyUs+iImI24NXtQ5XVXXvIXRvFnfXrnjGnjmtAwdf97P1wAl83v3XcR
hczTKnU+CjXlLuXeDWGTvo+cc++R9eNnR/tvmoZFujkTclNIl+gevcRMlQauHg47
VOAcCQuqi8PmBlfSCPDxSHr2sSVyPXZpI+M6dQ5dtHNN+Puy0w430wloQ4EHC0A4
mfdf30vJjoCDx/UJftU9ddMPGj+wu8+4hkogbxRIDrZl3ScA4SNKGnrKv91KM2jy
EotliJEv19A/YSy7+3xmWC0u4FSuTuS7N5xCFJ9C7prH/o9XAS+JyUwNuClMxrf0
+yVHXmv/ajRZ8asWZf0NXW/TOSShJF1GqPS3V/uuKiynPtwH2ToYZ8x9jNrhBsMD
8348nUTWPqLyuxCRRk530IiIpvOp7TShg7rYk5zd6eyxUl1rU4R5U9GTdajXN7zi
rqIJPsAns1RDXvExPnX1X5gJ31fD7LAUEnEd67oWtk4U3MboTqlKlN2NjD40j3GG
kggQG0KCNx3zfl0AGav6KyTDzPlplo+rZICSeMbVEFfkj83qFJGHA/iWwUnxcQfm
dya6Pr/rKr1vUKsiKyIsyjP7FcJv2SN0jV5I/46FPntkyWvVrvB4aNxP5gzOe57V
ubSpV2kEhqRt6cR3c7mdmNoKgWCMS8iUOs951t8OMLiiUMwqst4OQjBVhMKNPBpw
+OANyOXsDFe7iNx5NSkfDGhuKOutcjY4KXeW27qbU0AtWi/NC8tcUhiUuCwnh7Vo
AM94BVuigNLJRl1jCLmfOYc+wkCMA3Afg/Ke3C/Xi+CdAj7NSZgzqEAXcJh+Fgnn
nxhYCnI7648G4lGt6Nu8CAJY4GVRL8Z2RsLEboK7Yu0K6LQmwofoqz3soJ8fHu8h
O3mRaWPqqDEMh1IS7qtSBFFmZ0VL015bhj/rerCywL6KxXVfPe+gz/oEraWrOem3
nWb+R4NFp2AHfi0w2GF19e8eIxm6wf7ucg9fu0noICDy3cvxG5hmSi2iKW3bMuja
v0rZ9cAO8DbfzhW9frkDDK5LFMzcHR0oYSibtIYwdkVslQ6Sgzib9WbsOyLtIury
MC+5Hv0X5LAIUio76WpeHejgeYO84hewnUsp5LpxKDEcI8A727Ysdxoz2q2mp42K
6nLjNp35L5BxxRpJxaN7kSEY57iWjhva9i9Kw5RK/iC+mJQVLxiR40VsTSDt7XfN
UhT6AKJZd7xDdzAJlmmmlqDKtIa1qMtCMK2eF81r7zmelpVBQiWuT75kiIATL3dc
qXz+4R/kwat6Un9XLaVS52pUmWgt+YNtsgdQ93a8WVnj9DmPe26m2eMOyjaV2TGY
Pv0MJjNs9VU2w6HZt2gEsjbdB6SANmLR7D2ISSQUb+azia5TosUxG6HL0JGHXNV4
Gu2RbC4M95O8LhilUvivnbKJdsyvLS8EcMIE/guJkkaMNNZfiJgz6nVxF4NgivAS
QNo/t9nvnjdoJIBSkauwxqmGRELNTFnti4vC3ObOegQcuNKfa0usdkXFsTX87j3p
GJhljdiz7XgGGE18E1b8O0t3W9bO42uaKDQjFpQT92ibSVvewIePxd6GmWhJAIPU
RTjxyts1yco3rR5sXkxRX4FKuuxCX32zYvKanPPulIOh0B3MMrhyTcmGx7Yc62Zp
QIaOMprnbW97xxcsG7mn7RIVpCc0CIe+ObaAFP25+6Bzhrq6m7kh3j5E734Bd0ZE
biMIfVtECMX6ddDn+exmLyeAmkT9Riop0Dfg9H0bPBCQWyNs/eVFHP/VmynDjl0T
HC5O+c3xKHtK/BSMLw62HmSwcn8GOv/bxoyaD+JLEyy62fZmVTOf3guQ9WJewdZJ
NxQv6V6lEFP+m0Kv7izs1k6ZG5njJ7wZU4H5sDZCgR/z2XMBYdlflKSC2mkYYChK
Wqcx5Dh33aPXrhhfvVViP6fSenwtWqoX41oE3U4vy2RXeByqZZsln9VUkHsN4JMB
RvJPdfSMc93kqBz+B/gS2KxWbndyoZUEnyqTjlUIlwsH3kauQi4HkvVCzfA0C1AE
5maXAx8wXWi2p2fq4zY767C8mYTyUKa4+eP6YQOZsv7JtleCU1iuQuIv+mdKAJ1m
Pwx/95AGZ7W6Wq9eR4ifhW8GM5tldU4x3l6yuT624ZBRBHlRM4YTS90yubEGfZZS
X6CYOsCwLCaGFUlxG71Z3GGyVbnsjekZJ3W/NXfzQbKjS4meKm+yHIPxlOYGimEM
jqbxc1Mh/MK9CpleHkA9diWLbAFhj76yLcWwBntxbJrl+9zC4oIQ5N1ao/M93KBU
mNKCnzLoWrm06jStTPPwppX6uzEXjqrZX1sI25D6RDU2RgFtx/lg0s1Ia+zhN2rv
ZipBSBylbVPovZ4r7A5AIt5iyp68PMDGJgA2TOAy37r4w80BI1t4lTerZPG37ewe
+r3Fo4Tz/TKWXMqw2XdFmyjd465pgoMydZqiP1dWepG9rAznNrTCiccTB+F95o6Z
8+fPkxhp56v7WqzBsKaxrHBZ9YH+VGabk1rjpWiwnfjI19peVXNrYHLHr86w1W+S
GfjVwSMKt9N6/1QP7Qb69d+mzgQajtNofp0/vegtSOjwZV1rsJi/i5llwDYCnove
rzB9HlzPIBUyeogtqRTAWs20VUgeLADyJVHgTIllRDZ6I0SfJCf7RJRbnvJXsRmP
vgA8ge/Z6UBzBBMaAAv7zc1LdMSvNzNoOkAI3RoePpzjbKL6dkaP10Id43DO7/kY
M6L9GjvnAc2OomeMPLgIObilOr7/h7fJGn71OJO5ITSShKOBR546qAKluJADom9k
c48Iv6Em6PhL7NjvEIdfMbnPXpKhd1UM5Pdc6TxX0cl63Os6Y5C3wcXKNCaEoL4i
MhurK9E2HlwuJLBbkkdwq3xTKByUCz25gtoLFONbK5z+sHV5rzyndROlON/27VB9
+sAZ+tQkwBfTDVeg+H1tzS1MiLAdfNR1o8J7r8H2eISfSx1bZlGAKVBOuSWJPvsL
dJ/4T/v6YmnEeaL9m+oTIzrBpqvcP/9k7Sow73XHVq2aohrmkUyq7PO2yMDilq3Q
fu+mkwaIHFbroh166/DOPp9zJj6MONRwWJlReISU8cwKAclBVSW6W+LA7vpKvYHS
3ZU0eV2mM/DaKNX5Ko76P3HhuhopCUYb5eN8gTRThQZ4kT0zW1s5mm26mSKZa8Fa
T8hDa3qCbLNf33jR9e2ma0IRO6Xm/lnEIespitF/jHgw0sEDTnMYzSe5JRwP/GE9
sehauZaTASTx+ALslkdFIPvq0lqqDjStyuw46cNR5rreBE0rOXi6xKV77CcXTAvu
5rtYq7Uu0Icg+9JLeav1YElhmKbvk1eLo4kNR3bxjv2tA+xOYe+ocZKiAdyv6tYM
o7f+2itLZ2Fv32rmOmBfTSppFA4P1XqI6bwrSdq4/d7/D1kSQi9VxF6jyysprN4E
8nqRtFL50ynNMB1FSDQ4i9mHXH0Q6blTKGefgsS+n1CEAOJQ0S+kPf2Wa+yXcPRk
SG9jmRurVoa4+HZLPospXPWc+210AvpGJjTwV9s1tZ8pAcmvGUtKisRtXviFw7Kz
/X5v9id5U+hgjxhKNpsX8qV8dVe67xEmVyqN7TqxvSGhhXNw3x4CxMFJ2FENkW1E
CRshvJ7Qqfja+tykiby7GN8Udc+XiD7AGG/CSWgCPmr44zz5wQXpfdibmCPquUj6
nN8ix8ypLKJIVR8U2Z/A7j8B5lzx5+WtpHBDJJ/UjSr7fJNorNiX1n5XSY+lSKyk
7iz97J8vcY1GvM+gfC0SkvZiVgP2gLM7cqowLEvpVT7pbiNpSNEOKlTSre7rKRub
lSb9n05o33o+87NVQ9M94/p0SjkEvWXd0fVl9pwRnH6+4+QZAh7m8SMN6kQ5bvwq
48Famda+PEUUGNMoTo0aXSRCzt8DyZXgbAQnvYRDXj7nVYWp0AMKl1TBxbLacqSE
MafjaP8reyUqORtOkOAfcxC1cKmUYo2uM9Y/NK34sNlwJvASjscbtISa93a4y1CA
/yt1BmXtTExxF189/yKU4RYlhGaJXLx6noY8UPattL/7Y7HPdXynUtemzB+k0g5a
MhlqlNL4Ije9UCMumUpgFTvIZ+6Xf7U8ATmkNvcV7u02e8uk/qcGa0B5B4zuQ3Rg
geHurF0QLlCquzSbLXKqNFnHmoAmuxJ16DYVhuC05Jc3H4U8zJnbJ51YfL8fnmjx
M227BHPD9sFrx4uQTGBxmLUmjkBS1q+wZXW5Xv4Tqkr1ndtnvmCcud/RgaksVA3b
3WAa5jonHuh595HLn4Cl8/3EtiYhmkfx7zkIbFXd2eOuq4hu4/MOveVJIIPxeOoJ
3XfaTbbZEk8VNxe8BySTr8t3EmRkrhCkZLPqzFufsw+wN4rXquovEiejXwmWDK8V
DZ79EXwvjWF4cAV0AId7H8QXAH1mZjO1z/ikig0DKybu5U7I9Dh/1j51Y42Eadzf
RWR3Es3RoxNlTd8h/kJ788c4sMJVteUGwGo4mG55P9zj2/ZMsx1zMJ7ef2aOVXbn
qidaAW3II4HM6mleYpjzp14VnrdQiWX/DMYBFH+if/V6Wp3azLUR1uuXwpRH5ut8
Q99MQ08Ps894Sa7CoakFRcrqRzRqZKaVHojTkb8T6AiNVH+WnJlSV+5j2qcmNyLr
xt+/Kx9OZV+Ajx1mO54x7Mj3WiyqXkStXW2H5ccVHHQpyWHYVu5jIH8AMCmwdJ1X
fJ3IADViuwGRYfwTW/BZpz6V1dyJJex2ffr7OFOK/PvUZfc9vD4opI4XY+qYh8Ai
M68NmivhLWxfts3+3T6mYqIy2cTyg6pCcqLSzpy2k5gMyse6zZxCAg5EjCPQIftP
XCjJdM87AIQvBgzYoar+O4EQayyHfUgS4rOPdNlnS1h9ffdmAruVFvpdoHGfkYyA
o4m5nzFndwNRll2+89mZ2nPgoH5nVEtvBXMU4Dsq0P9xmROjt3Q3k4Hkwq2a6VAe
oP67klaGOq941c4P7a0QmPqaAHik0/GKKfO3InyImTYqFXebeO2oHMdZ01V1Fu1c
OD8yR1NXC/TamE8c2iR6hG4yg9Nwn9cv/LSjPSocj4OE+U0BDRk6q+ZQLhr59MLr
ot1rUr8lNHsE3gVKV88Kdftfrt4wXCOmKKkjCgwUp5z/q9lxs+Zt3knYLGobFM6D
gJeRwqUfTxdus7D2h2ZnquMeC5pxIV4Cie1oMzbN5fbyHNiJOezEVyZGyq524QyD
WryrMGfflTwUBI8QxplqQw/Y52nIJueziGuEUwCVlw66rgglePrrS3om9enws13d
DPadwjFqx/lSUNRL6wply2orgtJgTsGbLbr9YYiplZktyi3fpWEur67z5I7tIvyQ
xOJz1DtAvKmOtQFngGrWb/fA/PZmz8dROdgvUT+vFvJb5zmYVSSFDW7YdKREX2/V
u8rmfV2CusyGhnKg8vUstD3hN2AMOYFiPk5mxNw977JYCnxTEt2XHsF1/4G1mqtK
t8yXJidPwDc/KVEV+Mxh8+mzezA/3TVPZ1kYHNUvPkLrak67yDMg2XuNsKOKeZqd
5WW6VVfR3h4OFyB5/k5H/6ei8h0kfrFf6oyRHRuneyAeA29qKJn9kt8JJ40/xkgf
puE71PxI85MiVcsjej2nVRWIQwQD7+Cgh644iN4RpovhCD/uqQWNMtvpQn4RQyqb
iMX8ztQnSLFokdDaphGk7jQQqrj6t+X3NXfwrQ+EVO1MlKe8+yOCFysdLty1Oub2
Z9p7q33wIJ0BColOaszL+SmkqBgBy/a0ir1QXD8X1vKv1dcFR1xMbqVpo1zD5sDl
PZ/dTGq788qyTRCP1wiKxGr3u/tFubyA3jahCc4PpY8bqq1fUgMpaNAF3mguA2Rh
ZJbyp3XoIb7B4Vv9GfxE2EDNoC74/Bjh29BrpfZMBJ0lJC96aU3OTUqdjg5LSTT0
M5p8/VIHuNgreSi74wpzGAvanMEWT24QopPzYGvh+IQjRgQWCUZBstBmheixYrbv
AdMNfPUN8OFdRirBnS1ND+g7wrD1sB3L7iU+Lr7qlYqAcsE8muI0pqHP9Vw8Q4ZA
LTweHcsEDX6DEiSiTStAyVJ4zIBYcpGWNrQiRMxEwOsaX+CkXKNbsOR+cGXNorsH
GFTpc3BxIN1Fs6wm5ZsgO2nApjjddeW7IJb8faJW/BGy5RVY48SJtEDV9smC+X8X
MHqkloDuC72a+4A+KiEJfn3UnoW7j5xHwvnEkQt8PVPSZS2s94xLTOnU8XxPb5Sg
VQnSrA6aJwOVjN5OKb+2icl+PDeCKT4Y/gvK71xLWwWxGdrnHx58S+7+qSRMuwJf
OcsvRPbJ7FUPDeFOl4V9FfA4Wcd5qzyunSy8GUaumjuj2y+r39Rzb5xVz/YE4oXF
sWd7a5y2dbIbY7U4fb3C37i3L8lNsPZ5qKOdxJR1lcQv3Q7CLCZW9LiHVa650Ryt
SiRHwTJOJ2OmaCLDQszmcPWOsUxTtxLA9U0w6v2RyU0hDPmTDgIRCP7vHYx1MXWv
+g/ft3Bt07dB0NYQy8mEWY7TYoPdWilw1ZGbEc7cXrAOm4JyFpdiA1M8tyTtLLPS
RhYm8paO6HP93ZBexWuISIfZRCPMDxG1TP/bYW+/bs4CK7lCNtTclO1rJU36syqb
3IXVBivqSNMiC6+W0sX1/Vudh9UXhx4APhczFx31MvzYDtcQth+8gXLCGQHX9Iks
k12uHH9oRAHukV4eLz1Y7rEGJsNJSwY57imw+pMPq8GtplwoBWTzbn3mZx7jlDrR
FAPUjAg2lCT+NSn6kYEuT3VVBfArNhOIq0KQ1KCDn1aXmiFp6WitcKS8bOwHQuCC
nYAJfrVL15rd4w1Rd8Eq+Q7VdoAb8Hd1sLM1xfc66flHShNyeLfDbKgJXm42bI7H
C+m1L00UDS19oy7oihWk06OZcy8SgOBO+Dh7PUmLrOc8nbL93YcMXvOFYmdgnunO
Z8ko01SQ5EdHC0G1ZvqOJI7sOE0C3B2N+6cKH4ZAajQh+arz0bTwrIoTKnJ4XF1s
n26mzsVYIhaodNj4wDKv/+jwhesNnPReOUzy55kq46b7xM1/4GmLN6+YTj/jARlw
h9bV9arT/ja6XhA4nHrjA9C1jnrcksR66RGl/WIc6g/QmQRFOnp2NdYfA1k6t+S3
lEJXv5GuEUgikrAkSgKJK3316/eyYwv1eC92b2szHh9wUJ9zprLzf03s3FW/ZIXi
WiACdaG3hWHp9ivuR+UC85my2y9o//SHpFXWk/CiHcn/xu0lS9Zo3yZWnCdhE/fm
7fi6TqOvOTVlV9nkogsz+suBOALG51J3rfmWUe5QGMzGUEBmXzu/oamK3YvJxYvw
v7iN4SvBF4v6iweiXU+VG4vJUYo/W0kmQlA2kwKAx4K1EMjqv2MyXebwRILZAYtz
/j7/7N4AyhpFDt/vQYbCaWlU1CqHPQuHnA69gB4+yv/CNVwcC+ebD6jEjKDXNyMy
hbmSEMexIz1o4WT/PhaOE9ytJ/g9JW4P9sNCp5fzU11UKiJ8X2fpXVlo/P+3+iy5
uYEYYf6+CrHiiNdzwLs1QRmiZPvdtZcjLtT0Pecm8MBBAbPaV/t0X/tJrnlzLIp3
eDgtaNkSBPWQn5z3COndG0FW/E1oybhZvxue4mXttOY8Jxc+SPedAHY5RB4cpSLT
16kHhxewJLF+R+JApklKIPNMTr7rPT/SZMn3QqKlb9XnsvOtcvM2j+2xGWSPrlhh
ib1uRavS2FQWElszUfgnDkFoPB3RPS7wDexj0kX46uDCD2yfhL1qQdfJpNWjtJD+
E2UdkABAmUzLxz7POdimoHa5H7XItWGeJq+BuDOY5XaO/ldz3pMyHg0UAxX9xj/r
5SrDu1HeZRaAllUhZiy0tLBP8nVZaLLubGcwOXgbZqyUMVR4Kr8T3mduPAauOSoM
Mh3hme+c/+ABZqDRZhepVEnbqxcVkBo6yPjzwiUEYKeqjt5NAk+922CeSF16TURu
+P4Qb/BUUQY2awZeWUGTdwbbJyszS5wZ4yIHFn17WynWglp4WNcIyZCQmUHuXzjH
pPT7zIQzzO/VGEVjjcdUV0S4sRGALgHyCpqabNGlZlHIl/d5ym18XYZI2P87WDQK
FfEmFu6023VO7hYqwOvKluqXyr0yCY7CEp3dAhBol3gVVpYXpFCR1NnAPPI2Iwey
BlJxwx4mk+arRNro+TGUcWWANBLm1P3LLyTtnWBP/a0mlzX3JlTSPWCHqrv3jFfH
SFkAvGm7VXgI7UWFuD0qoXVsfE9818b1mik3pQdU+2ejGja/7Yxkbv6F4yo/JQ/T
8VtNQxBMtiAfKTHv4wjftHmG/MfGOlJttupCODPWJ+4QUd4W6aQhmvMZ12pUnlro
Cq3BZC2G4K5NyIlw7oTY3SUlQqA3+A+UnJEP5DxY499noGT2sXpD7j8ggpb4Jpmr
5wgo60aTB7rMjeLsM7aNHFixnQs/w4hfQ4YP4LafmEJueCmDMaBzyNq+vH0T83Nx
+UaxgInDX964ATV3VqdbizoG3CdmZ71wAeQuzBE5WCgL3nyovjH00C+mIefyIZ4f
29inItkNvEqwJjoTASQU1AEPW06Joe8TiMXHIHsT4Uwu9uwchXsqgEkT6XVmOyle
62gtTW23EV+MuFsdq3yqyV+A2P4Vk8mhsl7LU3ajuQaSuvdxsDF5v0n97ZXncubQ
r/frj1Wqf/qaJPFMy8nySofke3Ymu9e4bvH5tM/SXqiioip+42kBCSGL02Nnju7S
UhzTy3wLfZvgkdUaTilvWbQYCBFAwSgweffJ/qS2IBx5vNpS7DXCMzyxFthIHVLZ
khAB26rHz75QQ0lxHePaSa2QWrCgImQWkIMJR67mTHgWMAH4vQG3OdpY/bd9+LKY
9vUnjHfOned4wrkaeKTC+GdAMuU/+7O81GogXXi0d6lrhD6/uYywqjUI/O9DhF0J
bF5MDTO431e4A1whR8cO0i7Y1mIGIqQjITkJSXcrlsFy/35ab478Q0MzRuVr4ptr
9EKYL8tcIbdN4b6eo9VvtifgHHjo4rjl+FmW8q+NNSflD5Dgyeh5j7s6cmZ0mL4x
srNti6ICxrndT7rju2sIt82jfRV1fhxrQb9YnkI8NRJlDiz06ia6lfKsbSvfLU3u
qGq6MghNnWKleQ6y5ZQ1T+KtZNWV9+iKvDOy4BnSa2z4gopq5ZiOQxkQ2sDp/rMX
nCjmt6KLnqib5s3beEatLSB4JL+hxOPFCm0seJB39uVG+x/1m3AAcJGRd3nzFapN
2sQQ14hcPqiNI8EtvvS5jB8g9rTN+lCH8iHnu50s8x5+nDW2nMW34j/zBAXXLoN6
ONstE1hrqkrQcHyn/26R04eZ8ZiOateEG/fEXicUUKyZ6V5SvtAKS2+D5YroFv11
D5RAyeI17pb4OyedUX+25rwhFDt97jxwZaVREA3175tI6iOOshy23clHcCeI5PLE
fZ1WFGNkWWJ7WgOBPsgK+GRNX3nKUTTd5+UPXiJ2GcnOnFU1eBl0NvObw/PxbVVt
mPVlLJMRINGFBIRVqXs3Vo/6/A4b2evHVRYVrcQqjQsWiquolwuI2kxjq5Wd41Ct
ef4GVd754Lni3md/s2Nf9S75Xbq1DxqOQUGMguqpL4r4ytpk7nF2bUalUiTPYgKA
zWM0tXfOYzPZvyR2I1MQ/KeYRPMPZjAqLP49ESjZtJugRUU2nQlNaw+g7jIMz36A
4rAJmJV3/jm7iLA9ID5e/seoslCfcL0bkshgxvKsf3yU5q1xZqeyHz9PUuiaTbK+
FygvY+bbxE1KwidlwKJqP/Zi17rbPIVGKQhKFO2KzImHika712Jajd7qQqzjZZJY
X5Bb73ceJhn8Pn221f8XtEo5Ab8mEZbWaU6eV7nq4ouEZCiyIbIadzluXHdMWbTF
cHd9gLt0Xcv1FpcC7kgZkgaL8TbtTZkdk7NZdJRz1CNfl+BrqiuBaEVbgviWY901
hVTA+FyIOshvVVe+KDOqM+yjoQigGBXhUOJsW1MUuktqB52RZ3wi7qHw1ePVgSBa
TWEULsDhYVBnIui4E440tqqgwhtZ7I7nXkv8lwFNn6grTrqIdWZOWAvbN6FKmvpI
IGfIVEJxhst4/GpT0F66GP3sCWOPmPOPYZfGw5TgYMeCEYJpSl1jTJyOh4bVGdZW
kpfZDGmAeT9wUccdrZbtqQ+n13D+U4/3SnX1xc1NM5p0ogc5+qRXSph0dOvK6Uy9
Pzmg3kieH3/Kc/s66YJQxi5c5Td39qgCd3Wb+c3CCKYG4aYkxc4u8x84aFEJ/Quc
/3MFtfaAPxP23E0yLcgbixMgpf+FuNUIBXL54DIFa6aKsJRP57bliTBFdV2JUYHr
M9AKQhosXCslGz42ha/PyOmJJ+OOHArhAX7V1AY9QaVSrWBSVY0hSzNDrHrLq6f3
wogRQgLG9PfNTQplY14THMheivQ/MhnYT5cYh6xFA9/CESHek+bEB09Fnw/+79RI
drPaFmpviME6tv2Iqp0NUD7cECiyuJ8A6ED/fzzz7Ld4XzmG4P2nLcGjkNyHc2PL
SbK4/jNG8aXAFWBPDN3FHzAVhEGf1u+8vnUOnoxRMaDt4TM36Z1IkjnahTDCTkjJ
fca9GdAIvHqUqqpi4egnpVTPt3feRV3xil36yYxzv1RbKGROAkQWzJPxZTNX9p32
aMRtzy/gzRbTW73HOPyGjtI2rEiGlgHhscqi12GFU840uyr9hIc1NgemvUcQLPYW
jqVXyj0PufhiL9VL8q8U+o4g15oLMKwEmEoV5R7E25c53LL2RHEYTRCPKV8xqACH
rEKnPoSLC0rtMZ8fXtKSyscR1B3w7KgjsXBHtiMu7+7bPLm47k6F2mo9BC2HU+d0
bgIEKe62kCKfik3m413+TIx+eejxnsybxC1ir2HZlGVOqPL5wUZQTaYcg8DPVXvr
HRKQg7mcLPojvBsMVbfp9d9BLGsWU8ejzpfbYpgx9Sbc8Swnesq+iUTPZcDPIyoN
ke0Eouw2TqSNmPor6vj20VbZHa8XK8eV/KzP1bt1r/+CXHsezAyga52vQyQKSMhY
W3N8qKoZf8jx0OAhXhSKfJKwGmhKuqAi7VmIzej5dQsYRUUH7J0UX0QEyBqbLlM8
xJdoLXR/9BvVqNSH8OnQrVSBWEATLyjRiU630nQJpCzD7g41ZzmP7W04qHNPuVFW
CW5Rjb8TC+lMDYWOQZhhfJOaXHM/kaXDau82PYsK3zLISkSwPP+ec+YtPlllQDtW
oBL0NA8gbL8BC1SxCPJb/MRXtSrVa6UMGLPf+obH3uZLrnl8SgVlCLxgauwIYj8O
gxvtjvmlGKIyqvR36oBJirTpQQfBw56R7J7wjgwshuCJOQm4w5ot6cVrm3w5ezIa
HS9ttDlw9xJSQZEFyAqWUf162g3x5Dq64gH0aN1WRNiACpG+kBwr9Md1A55oawkv
o2PRQeNIs2ytkc10nWNvDXqK0eeuEJS4NxXO6zD8Q9vPeNXPRvRfOpU4NIMitz5r
Q4/naIgOdtS9yQbkWyHglEmvtC2JV9LCpEfV/phCNj+CwKrgKSRjg2iAf+9vvRiX
zSmIl0Y/hyqzvLJ6dprTPs4Wzi3BRrvYuhsaAJhvL8Vhq5SFB/JsvWx0JC/TkkAR
1McOY9MxmaiwjFNEGAE56vi/F22mGXWMkqQdB9hU0/v5O/8UJA4AWa9SfjeCMOsw
ijoSWQ1OyFh9Np9sI90tpVjgXhPqq3NOXjiOqRmIhW0SIZFI1hcsP5pnITzOjYkh
QWivuhENKqUrBg5+24bpTuYv+WJbK2kmeWZiI6zYQchDsYAxv6RudHFrSxUfURVk
HyytP66uWQTl1/f4etdtktT8qW4qQy/LrCdvFAcAWYTG23w2/BjbznULH7dNRyET
31NpHDotyzaHJT2YLMQyyjVwLKxGrHLHJoqNoKeaqQtOkh/VlNQHuXPIZf1A3Ap1
xoaZgixU/dM/KAkErxCdWGzctbqw97fLGBRyI+/DXK/bEphDRKbScZNfNZhE7a4Y
b8IfbcwrH6Sa7hLnYiQwAPBlvdkC9HO/T6/dbEOZnH2VQnpMREqNbk/ezBOsHnAo
1EDGu+BYIHsAveofmDxsVJQJ3tokZgcRhTeo46W6dI9SKIXrMF2vpwbCHHsLN00+
Sp/rBbqZMsR1mgcvAS8ybDuV1ABicD+21pgNTueEDi7OQLJk8zX63XN3eNeirvdJ
lpInnmk4SAgcyDgB1zFQiXohjUPiGl2PuMxctzCwMUT6zIxAEUHWDg0amOvQhCBz
jsDWRCkVmdG6D3icfS+TWNxKq9Ty1ACYg8z6a1ARmmidc6rf4NMtkm7Vr0LcVGTD
2e39ErlVbCtHHYLlAuWx6DpvATfPfs7CRw+z3oD8JIop3AMwPg/jo4SMDJzhzpvN
rvPajqzsyPdXv5RYdHaHi6V+oM2NOztUahJSXkjkdunSe6Swwed62pd/2Xyn3UQJ
a2Am1jIWaqi7KPdBjfh6xICGf2d9wekq/1QzF6/bkRTtiHKltQ4MVT2FSv+JbZBD
YwjZM8Gn9z+Ibv8gm8nQKHP2ZOGj/NWDKAsAGG7goYA6HJpfKuJw3EdaxqXHUbya
aT9IH4Ym3nYIowzuO56GjO+FK7S66l+RkybAcSJpwASN491R6tgOwTWfpElYZiBQ
woxyJK+3sRd9k92rFKqlZnyBQaVezPKinrzXKF7jDQwuA9NQORE6IlvKzyjO1viW
/etwaxqidRzzmbVUwrGrhAwyD9szJlguwWSqcdi9fbXwMNeybVMoeCa8+DCTwUV1
rZ7DWOStIWva1IV5Jc2XY6zLjnpMav9S1YNHsU9MTpFIMCRA80cDO89V8Yfmn9VK
F4KEXqvfbnkV8NNDMnnv0CfLm1gduaj5ARzkt/YSJxrVbA6EoTf+43hclQIY6gME
53ZcS7tkfvMLu2r5mbJcirVUQlwUj7WWfwIUhCsOeMIN+ZPC0OJyXV0M3j848yMR
uiSkUfJVZg9BzaqItVGxr+reP49O9OzBc8gEiPtArAGtQvKt/+fsZOxBsOP5Zyae
IqkCHglmxnXNgtpMTrYdZH/nPFL+r7kKy6Tfkigwir2yFeimiETUUjB1jvjbp5au
xX9Mh9n3ectTgAdanW6JU1ONcXulpUaq+3Uk/KmA8Dy7DO1YKw04hI8mGoA6u0qI
D+7J5UqaehFgeQlcde1G9RrWg4hjccKsQp3z6E/rNIZvuEwauW3erpMggZICMrnZ
bVTylQtGCulJ+JEJDbPi/nHuZmhiMIeCd54UEVjEViX3SmqjLbFwaoAjQA9CCOSu
DL+SKw6wW/KOr9DnMEFPe+ZoXiwTQjE0Jh9aMgI2jvAW+wpNv+48lpYS7P9ZWdHr
heh1KdNli9UaPUntaiPCie6oQzFkB5rgqRfdwzYGaHZULkmko61swkvsgX0x4tOr
zPAYRLxxmhCw6nUXO3XqHN6H3LHJMCIT3dPkhOrS11EaUpad3cski48kxePCimlt
hc+XPzmrW+RdiyPHtHTVs31/jujMDcLjUhzycGk8FpDv4Em6WKjWyZ/1xznNxDEy
zvaF0cD33O5HmHGlLRsc9amPSesvkD32tWtyz9K3KUF7jzes05TdpVLyzCk6shH6
1h0beIkIAfh3bY9487xV0QrkI61VjjfilLM52n6ZSZ3qxfGHiRlzmPF/a4cJXixL
SU3ZsUseamCYHINP82uRe3B6vc9sM7l2h9jFZgtXX91IyP6zJLeN1r5NgINCZIdZ
kaAncKja+SVyDkgTqEZgKUbMEMWSJ5zFT1bOyx7Xb+Ih+wljOTQW+jkWPjPkJd5H
K14L0xYWHXK/SRotqf3o2N/c8KtJYt6ij1WzSHAc8rtA37fU8lwvQM+Cu1k5OoXo
Ilx3AspYP5AeOse5yb5V4TCv7bUwD0BFL16C0Qu4gWtMlX4jDOMMKJ7O154ihey9
KxfrdwVlZYLG9SMrTYvi1HzC8++wbSJBmEtYORFBBaSsiJaWWXfD2rirEfPZ3+b5
MDi8AIdz/hvLtTj0rJIk2EZmvSHeWg0fW+1WwIrRIU8QOXCeIB8m5AKx24w9DwTs
j+HdZNvQj4336/ZLcCar2oQ+oDD5FdoC1Nf4EaImCSqUnht9XzXrv58qJuBRsWq7
tPRG1jo+DjpbIa9iHOfh/nMkOvwhjvSBbPy+NOPZWc6iyF4+rBNhtxcsgCV7bDdJ
NvJd/aWkfpx80B1Xgw8uJH9mUct2XJgpgXsS51ng0LmKsqPEGc4VZPEedMEVdnqD
eiyYav1QnGCNycJTYlcqMrtR9ucUa/aYwKSjCo/3jRx5z0imqrVzm0LuUAoxX2/N
BnCW34IpCPu0a3AHqQDhdgpcnjtZzJ2aW62xcpJBz73ObaRAI2rhbUl4RsBIOYFV
UsPbCSwFMgyixA1YGMx649ojIoPdrkh4gRuZ1LbfK3ISZ25cAvGBLdJMASbqzSAp
2sVOL++r4BVOrAIkYnaksvHiG0pm7+WV1CJ4XUQOMl9jQbbpDv46lAxQ7wf5Kgq7
rV3CC55gnWCJe/SUWgIb64Ou2AVWj3UZrCwucanUM0uKCxCDBsQLLpFWmmSVCCwT
FcCJOvFocWO/JI+U2Q/ZkbBxN+v1alNgdaIMzDe9RdXDmXNybsfg5mF/YEs0Xc8l
xN8bwpBw32NGKjyizK268YEAbBxm6eWE0As5/ULh06j8DcNt94XEuI43qPH6mXeA
oDQDC+uYeoFByiqLn5Go8a1ZHB8Z0D7zeG6lNTeYookPMz++g0ty9nPlfVHb7dnq
AWeZ66ULrOTBgynWdEXaDLuFfYLqspVGZwWpNm4BEmjTuY6TBjENj288piHrLBGm
RjawsRthxlJchYzOEKy9K+EPdt1gabDezgci7PeeB5SvHMGg1PYa7p211pI+Tm6z
xn9bjFIZBzXMT8DqXqzj9dJDXkwx7HgCiNsEvl9ZfDlSqur3rd2oA7A7nckLDJhB
WsqWvqfaLArcWAjuQFi3xD6pXCeZCUSPu6TFKCCxIvL3ClE2+pLad3wrXmbn4QAI
rc9rh+D86h52Kxjr6SfYBg9B1hJZ8z4z8blWoYqUxGFHgHftqjI0oHC95PoURBMt
mIuHKh1fmgBdnRDJZSxP4UiR/NFCWplABxUzuka1jPDw79ngKNNfUxFvvTuwjV3F
wtC2EFiyYoVnkUswY1nYN3hsDVy1EJDufouIDNhw+7TXtMmKXn3bAqjGEFgeMBb1
ZX1hMvCvz6h3/X34NS/hdxWCBpOiq3ZSXybW8uxN9lp/BRLnexOEY6UdQnx5kDrR
uxu+QHTiuQ6DJlrDWfDlaFGdz/PG7on9chrM6FPdkM7EyhwG1SMXK6iPVvABL3uA
7yUmXm5nBVnsTYVuTlMHLmQNqdz0l2E4oTloe632L9xDf4BI0ptIf3uRgmyGtooG
35I+Y6JmCzxMeZn+jYqxIzNAi2Tykocui1e0nhjXDeDf1OKwM3e5cr6qAU/4JIth
TrWSOn4/moq3SkllXuivnBEPy4m9KYX8sRj2mlTnObN+tOVqF5eoautVtTB7dy/Z
ORtFb6Oc90SnmxuikS5dofUpMY4lfzm0pZBsc2aMIVtJ8JnKxmemFU+zB39+KLT9
2KpquulEX2Q5YXZxfMZ/kM7VXjrKf6ib+nxeWoVKjED0uYV5cN1fbWaiLfcrv93I
aC90BtLAcW7q6o8IMZu6Kuikx29wN6vuJhaD9Mtpcgk1WldNVnzSI8+jj0g0dI94
SDmnLPawGZ53yAm4I6i1mS5yStrTWb7Cvv2TCw1M99howueGjB/WqmtWDbbkQ+LN
tF3i+Bl/Bl/NypqjOaB1gwcJEI9rA/pfpcDxlVzW4Ul85RcidCL8iotH1hu5zzwS
jvBvKENiy8qQqE8wJnys/NvhuN1ncTgX/y/o4/ymMXVdvqZTrZlUQfnIkUPE6aNP
MikBC/REbTRmnF+S3GrPL32OtE/cXQu/gazk/MUir8XHnj7qxDnsEoDN7JhUG9NB
Rj5Q5uZyOpanWTEGwtZkzxrEC8e5it9A5RDiyw5Dw9v0iYiCQsBQKu+Vy7kgzoVr
ELJMCEK27vpUwRaMOzid6naApBFJa0KQZAkJ/WD+mSrcXCQJGfobUGxgquI/q89v
cAONoQ1IKsqtGCjxDV7gsnH7c4+uNQUDNNImADOORvxlGUQvnQS7y2Kr11Nihzyc
Yf7iv6+DkXX7M9UK0H/81UlkWgokOnLJ12Y+oVFWQvGhpWP4T+ueyhVuL5n9j6Dk
8MZwDjUSNgozhX+qwRT4zIrirQAuGJN9B2la/0a5BH+GSqffJ4yw8Zo5g99yuef8
bqirXbD0sXdszEmjvaAaVH1seiJVy5szuz9+ojzykAg9MynaRxKeIjzDwPfEJRyi
shsRRH+T5147NC8pp+16uJ6mZ4jqk3maRuIuY26BwiWbLLu3rYTmoDaq0LA7HvjP
Kv5qo/I8fO8WoJI3Bz423JUzbueBDFZWpymMOVPSLj9UyzTYjyYNMShvB9Q1ajJG
oWDXAwnIPmPK6D8LWTrsUC2XeTigRYJGAifz4La3DU3zU34tEiuIrZtM7XxeYnqT
yof1uOPjrtH335da+T+RV8SeHDwrV8N+5OwnlLrGDwBokJErV0jbBVkygh0o5o65
MEn4wPMes++SsAh7y8cvlQAzL24apY6Gw7jURKwv2ZjIk9vfA00+Jy6Q64qxqTp/
iemwsdOLY8btwikVZxLSWa4KKhKqp357NfsoQX8aDboxYDRxHJN/zNmWlkkDh37f
b9Bd8ZUse3BpoCN0MJ57X0HqKBChsfsJT/bZ73ebwZmAdrLiGWVp5DP3ZeqDH0Gz
eHMelIHKkltZIuB1jt0kKDSr4EbtNaV1i2knbepPrjdkz3k+2xP1RMgG/fHvgt+j
uz5k9/Eki7S9uomoirAcwTOVIAPpM6+BgN+jCJtjEE2bLHQjQcgi3NioUqUN9tZf
sl9ogyDxbg54TeQ00PpoUyU5Q4dKZS6SYPnuKMPf1MGDQP9T806/j/3l0lbRmuUN
FoxftzWzDl8R6RKt1+/bAUGD35IeHdV5C8BYs0T99BziYXO4fimoP6IJzPdQYfhk
+8ZUxobOK/oYvYu7oklHl4mOGNjUrqdSpU1WTXO85JPqgPmXh+rlJdaovtVwrv6i
QXq04AZBxP8oYfBv+I7ZvVcmIGnSjwz5Nv1qIiX8Gufpv6dRAFbZCn+iG+MNUHzy
D3vteGyhGiX99tBWPCBVXn+8wXMxB5evDOuzskfHT7CuLLTdlmGLub9cCecHYiEO
hjqwF6ulB20PjDxZydwzscUSYpIs8ceAKAR6rRUt+W2+K29BptozD8q9yQ6rM004
yVzVcjnj9gkLqyCdI+dobLme9CZTPWQTvSYdQBquVH7av+nI6QVsBIQbwOahZG/Z
gOaiayBqk67+7r5TO5U1CTdIMWy3+hv4pNhc5sjlgPbCbenSIHVlM1OkH2y1DOCX
N1mq1b9/NGV9QGgjdvXT7zSRnWvk9yqrInCboQDJIgWTbRcSKHCmJM83nKTYK027
h3iImn8Gc+5Tl5XUX8TJ+RDsb1pePstoqIGDf9QIJyBtc6fgpV/q2So3xhIldIsL
q6hcEJ7Cwuxiz6w1DSmqOx9dcb6txQLoeG/0Mtah9ukNpvp0X4WlSfe/NeyHcGQa
s5299NmOD/ptw/XAEdlBwN2315UFjOwhakLh/iai5izoZoRqwF7v6sMWrwqE4buf
VCvyIMQzOfveTeDrjlXqF+nq5QiIb2apyoWZK99byf07df4vpqRoW8sSMTWwAJQX
xZqY3ssohY5tUy6+CztxNJbZcuePlWos/cjQ1G2rIN8Hwt0i03AqYDhcxOQWio9o
kDPxEczgByJtML+zVzIb0dNDMXNVqBfQut9+F2MWiygzQdO1QFdcDBz41FMrUjxn
kxYcbHzuquUqgwBl/pDyLac+vxesupQQkm1Hy832Cyq47XQ4Ley8iMthx/1yUAaO
dzQHSxA9QjR+eYaYAwdpp5e1l0voogq5xjBVtiw989OXqLtR3CYqifOwLLYmOmmC
uj0vAYnA+p6se7uiexTp3kiBsekU52xZ2s9rsrA82blnDYXxCNGpWdtcNvYlGQfr
0EYrURniMy3BN6tr+FccY0jGvdFBovO/eSAeRdTsXITOhftGvrw9y81c235vlNMI
c8CfxT4YsBKG7MMIiUQ9EXd/XV6dqi/S8kEqwcpvF0mMY8t3E3mf56mYaGPA2SJw
n7AX+98JttgHI299vO5aHjaqPNkAwitvgKNNdfGzOqUD1IAWODPsjhGnnpJJmQ/X
21O81JOaC+NcxKiSt/PE+2jNoiVl0f9Jh6sqZiJmUomdkMYhfRixWQplFtp+Zvt6
ZZBsQ7VHurgjIbJwtvEvyMRx0XOlWUctgkq9Oj/6En69tpOzTLca6mOm35GBMEBr
cLVxXl+P7dKpU67V3brW7nE+xlER7P1cceBnuMFt7W9daj2tyOHbhnV202+0cIPF
Q0sQJTTZSBbLxLACOLmOd7OaJsFPMVVSOLKgw2ujkWQxvkyJ1BaqGoA4nc99CTHN
h+HguPlWVTJlFzS8pLz1dlzhH84mtMVirn7P0Epy4IZnQr+5M7O/5N3JgmhvPxyo
+FSLwk/6B5P4Rg6PMV6yHjeoqUgNO2IW/p7Sg3T5QNLZpWJ75RSak89IyarWwW94
V+mqJDG6F998B3UqLiraRCGqTeHQDs1gdfkbTdIhsqkPEv+AIRaFVOI9SXtuqBAw
4AX8MK1ep4ONl6/Km2Urmn5vj1FAL8+d9tt87fneJaUXBNB5B40DWak5RAhnw0EU
5TQ5TBIxUFieyw+IZvWWFppHLX5sFnp/fnRXjB9P/S6auU9Wxu5kiw5Z9HW5VewC
xHD16uMFhyNrF64+sButB+XVanpkFTclvM/dKCfYR3n9WC5pvwXegDU5caCasBtk
R+IYO9iggl16fn8fULBTKv37xYjGhBn1lz3IBSLo3l/lzJOpr1r79hy1HxRoLoJR
Npgf4pj2sCBO13MXWaKCpku/RdaXUdOz84l3YAlOkSoDjWKqsJhovGnkDAUK3tSl
1+anI/I4AHHV34uMJCO7Irn1USSqyg0ayJnik5D8d2Y+K+EQwYTUbevUWQ5atHo0
bUzAWIh7EvlbtwjRlHKEI25+uBhezc4F5cofW5JL9HSNjijfnwvrz2Gu6ns2Z3qM
LcBXb1o8sFEG3MJuU2e+P42K/CeXyR4s0OiWJ6Y+8A1p+kOr0m/vsSQhFI9SILsp
AEkryxsnqUx0pfGtP4c8/AV//+ZC622mn5u/4KSAJvYKHUeDaqp6lPxYBFERFh0x
r9Jn9Vvq5iQpzsAmZBgSM2e3IEaDW+HsFS7XBLvrVO+GrsDimsSzMCRpp0SuNY8R
L7lERuPpWG3W0pgcFBz+gumplAxdHPYS5ipHSNQpRFwJFty7aFPlj14Y32Si4vi/
IgHsV4heiRwQnaQRZYKCJL1jXNMu7cxpshKuX7qqi2UdY+0Sq4eJ8kHj4VDRZ30F
BXjF9gTPVOuFdIfnNP86rDev8KBqcXZ1Q9fa8yfnIszN9HoSpb3IwMGyllo24Pe3
BcZvnnZRdU9xwcY+wvwPl5dr5ghTvVmttbj1Rx6/ejvz8Muo1ox5KfqdAjPw3X4H
wfocIB2QINWyppEog2fqnTTjWzG2Y7rsgim9CPq262TjTQj+N8jQGOO+HzdfRdCw
2Av/U2TBuGpBnTc2mCllUoarQSIe0kZub7bimJdFh1AktIQw4OAntK2pBmTofEty
T8YHY7Dayfx1m/UMWQmGnab3hTY9Y588qFErc0ghpb7egLntTiDJJhxigQvcQ+7u
Y37nivECTzcDBFY2SmXwL7ORddP2mvanuq2UPKkHj193bh14OCut8iICjBP1dNop
z4RVmTcXUj0hcMlUqr1/fTZ52UpXYv27fVOKsPR1Pyd2VpaJMQeEd6x3O3N3WuBa
C1Cn2YEtdQ8McYeRN3u5JBGhfcUsSyGZgcwUc+a+zAtZuuqzowDse5SpNY43tTeF
688UdujeNTS2mlr2inYRpltIIByTm3NejueeTCoHNN4DNJAnjX1MQpQoIHMPEecH
EVT36RNPwtbBoWpvhHQUe5Poipi5TJsgElpBugxPB+ZtAsJlWAeH6nzv7MeYYflA
mj28xgkE6D/4s77GrDfx8ZiV9QJSBHmaMqzali0X2trbXpjz6NGXS6257GW6AguS
w/Xx2zeaqqONjlt5sm6aWyJuVf/evmTeZx7Bcj0rnWWRBKFzxuhAAq270N8GqC6E
w2z5m+df/1ieZtx29kcoYbd4/YN/EehPpxYNGBZMiC9WmIlvTKxOp3NRn/PUfyNs
Nj2+ra243+Scfdzm2szUDgBR5L77Zjez4tRg1lD/ZOLJptfZHwUepUn1g32TAvEa
p4x2Z85XuW0YyVIqeT8JtYsmCMx10JukPdaFQNv/DcVX6WTsw9PsMKCvy6Xbp545
DRt5g5JMAV2wxCcvr8mjazuiydax2j5cWFSNoyvj8i8KaRtBBGpBvl5seOrAVCQq
ghTO/3NRKe1vXUwtLowdogs0gJDiMa2BFYCn7GttQKa3kzpcZN90FlwxHj5KXSh3
ohXCniaUyCtzDq01ODL2Pop6WwDXrpZrmmGVWwm8pBcLveErWg0PG15/WpfMEwqu
cI34EE13pDrNW2NQuNe37eNMfwzo2rLSNdeyC9zMYjHCQqCyfTV25f6tu6LD7UWa
AAtEqMNl3gtZ5kM8dDWAQdBxrjpSEr6RCicRSL/H/C3wC2qkSTRHLd5Ibs4yw2vN
/ABCGKhHgwpSZLvyxh9u5f+Fw581K+cJRCBIuZxHfwJjN8STcvRjRC/7YJKF/14e
1R3CJ4t7s6+nbxcTHibq9EIeYqcOIyCI436JUmYsLVzv4vmPqBrj8j6/AUUrckuT
sb2/hdLnliwX7Fgt3sfkIpS12/JFlk99eecZou/5B22UMJwuQUZYi27Zoacnpmwk
PZnunAEbiNb5oXUXJbFEuhWao/c8hW4TrRky2FNRCML9QAMHt4Ycn4oUebP6dINI
KgueD/X/FU94aFUfXIzwZiYTgjrFSFrJ25v39JdrzbfQe31ZEI/w2LF1d88FH4ol
EhjzzphF9T/WQgbIXDxyMqe1r/gNadsbqO3RcXyLRrVSH4VqU/1vD+85ArmOBmwa
5KeEmTV+JMyOtc+Y4e4ouvwHNe3I4ApN7hsOtiEojg3SYKO08kYtbkTqptqBx/eg
OH1qzod4stVHjFok7ZymDTpFWh+B6NcUYC9QbtTtpWsS3T9Fc5q1NG5+/QYQBQc3
+lF3nxHHivO0Z8lk3Mo2tj9jxSPmF3R+Y4OZync1F/catkcCBBU27ZJ35O02Klaj
vTFyuy7HgkK1sN8HhC2TjUZQyo2KfvbGaAG/tBE13XzO6at0R0kGVqxszz3DAuXI
kZjbA7QRDzIn6nY+Gf883dJZkoBB4Tq6di2XnfY2oafGXHbhPfb4e/A5O8UpQsu2
UscXvdjN4rYOAWvmDwZeNuItjlOOldjS/3U5O0vpBfhaGsX5SI0xEvOny+ka0mXH
WTpQ216l93A05tEvdN+BkBxqeVRpj9v4n8y4UnozNJKap6iE6Ad4ZpUGOF/rrp3A
7jsYvA+7PSk1paAq0XAyKK8LwEKrWnlmJCdLgyui+ypFeRroKhSMOD7gX/zDqSoN
tB/+dCyQWkLt/OgjoXnOuppjPPh1MXMChKKyzpsR60Tw/oJIJoVRcO8GM0ifMvtV
BjXzTog0uWDVMU9kwcCIjSVknY43DL7qGtLauEMoITn2M6j6XE7M7xBRAPVUYQHe
SgrI0h9es3ZS0VbI2cTnHB3bxCShB1z5H3YebnSdppzfxhlB4ivkzsAzCfKeh4H1
qunc1P2Q6e/i13uPe7Luu+twa6/P2r4gsc4lOiqVLFwgvQbP9oD60ttJksBflGzv
DojwyigwsIyLG3jAZF0oJWt2d+tRZEZ1ElDfDAfsY768myDqubD3cW5xtU2usmCd
pWzOWfNHqYjJtEwhLyQkr2C+VKaF3viIHzIcVP75qDXG1143vCOXKecmpOT1L5xd
7AG3vz3pegOj/YUYglVoQnYvPV6cM7T1EjvqOVcGjozTWYXmoG1gMc0E2CW0vGpP
LJl7ZAJkRnM9DIxuAw4vqfuPzm4E/BDNZz8BlTgNB7snd4OnandNR/YFJ0PJtO/c
EsdNQFvXeGH4ZxdHpnZc38tRQ+/lIVLCGna0bLuFkzj2l/7Vh+Bgk8C4rMPcwIrh
cqJocciGAnKUAhgv6BSA9eZ5Y6L5Nrh0RVY0ibeR1+jS5QLur3HO9xdigwK20E5g
qIJYpO9c+6XQoedsRbhpBxe0UBsc6m32hf1QigCgZFG6TgR/sZXzkPsu2QupBPQU
whbkEcVfscKvypxY6q8WCOx/KKkq+u6g0E3tfJZ2MOuVWIKvJ7aE/BD25l8zn0W3
W+g3JCtOPJPt3ZRhV8sUZWUmVgLUHaqNMGXZVJSOamyANpXS4r3Q3WvkBl+bRQ15
p/KUE3HDGrs7XO7D+u5ROrZMEswkimOQlaF/9AqE/dCmjgHWwEU9uIzbt9l/BJmh
ZCeVvCAdPObIdC4bzJHhXR+YkFs+uCSE3cfNw5d31FDMOiwLhzMVzce4kvr4X3pc
GzinYOqrDU868UAzPLr/8m1IZvTsn6JFKN+d2PcGg+FRE6hJ8xX3JBWlq8K6DbZc
qQZZO+hN7JtRMjSydHFcBWvx34gyuI7/MKeA6JR30eqz6CXu943/KirB33o9X0cY
kSCdDkLk45q7VGT3P79W+Ch2LXK9U7EAeGf4Vj9EeS2PyazcC4n/4d/MzBZJYUZf
XNTN/R/WHYnlvy+d1P1ihAMkerZlhylsxIdp+Ofb+bEDhOJx7QUOorVOvrPiAEyu
IHhhPapnfqIZ9dMvFKxvSziE+/Jn9/KgWcie6Nkl50EAua59TMArU19TD4ZC+TO3
kx6xeeTOfUQNi922OzeyRgcYInhbR2Kt1GNX3GDi8i58bxEubQtlZM2xz7RKpxgK
RZxblwYwbXrBRFFOC3TBXTUc8wf5GECxCH1sOJtQlXTGvLmtf32B/Vs8aHbFtlQp
zeBXUP4/CQCecrp92vssW3CaHRWAUNi2FziIdB4+i4HUS5eFH6Iymo8wIsez/T4t
GXS5y4PVcV1lr4AN5UwGuv4G+bO5BD7j1lV/JZ01geJgIrNtpgdfRbFiyrTceLdP
lKAEmA0iEbm5NSS3ubIbIuM13RoKdaif3v/WYxHSYmTVRamo1q7FSi+L2P3R3fSY
mx8Q3yAMFm+752qno53OoDFoepaLbnLOlLml8bJToI4ibEe0BBeD/XybPWISzU9v
lZDyaMQwvYhLm/ZWO11hW78I6ZKhm9AodLBwnCEZqneRBfBen//G9a5a08sFFmdq
2GjukTPsox6pPEwcjPJ4mbm7YqGNZXS643HHk8tDKBrnSx1fCtpE4qBE4OBBLLHA
88BlhbPqSdnPDX/4gg9DFqMysSr08eKOAs4kbEv7xgN428sVX3p1DGD4aeQSvYOW
FJMH51zhzTBPviUVFpYeo8XjEI7dyGHvVnr24mfCShBHnEmEX/IMaQBm14lgtLAO
/CgX2O/x9rvmqRkjYdgJ11aXhWAdBcZ/mImXIpdKKsjS94vEAFYV7ZewywZX+JJG
3P+uHkDUEYp9lu4CF4aDsodkvAZ4eSsphwDMC0LNVlikUXRACecpjPSxPdXDy0U+
7gYuPUL364wq9zbEuq4wbn1AaOefFgortZaBG7RSkkxHiDF1Ubj4iOrCoNTL1n12
3UJdCRo0oWdaMYd+8fHxf7Q3HvZruFNhsKVMggOIpJ05lh6u4T3D3CayWIUYYG6z
VQQ81hXhbsR54jNlLdvMhaYjIPhYc66lJCspFSTuWKNvHsZzVXeY1evEAMXfA9H5
E2Dof7MuODyp5RehS7ER7Uog9cRTngdIQJuRCP/0vCGvgS7ZG/KybDEZOFugDKUp
4+/+fx95yUAJKUFf7egpyvLCE660w8DC1DFp4wYu6msu4ogrGJcGU6Mf+ARGGO2Z
EJY2Ir3fOiImtJz13whgs2S1ibDZuIlevaw1Y1SeuHM7b50peZIM5M2xjb39l578
ib6/BVyJp63L8BHebwCothomqlcxLEvE8HizdtUPt0539VyE6rLntlMkCUJU3hZd
rU8PuAEA65NpRMkpl68/UQXyHVkWQDoOaWMrHNvp5VYRILsTIgKcLaU9UZQE2Aoe
/TdWrOcF8phR59O5u2WvJFrx8aMERQGPocIxysPQsWfX04AQmgF+2oGI6YEgON0d
KqzHmsB9/kfDuMSuIb2Ir/7fDw2WmD61cormAnsA/mh+z1GIHTGF6rUa3O1vVAOT
Ajte/4sqgXwsgok/Dl2PGSIoupU6OOQarKuUTlGog3JyQx/9azd5ddHjRRietDc2
/W+CGb71qV8l9bqYrmUtZmX4M6kwjnNtLz2BJiOMXI4JKTjnIQNVFQl3OHnP+omp
j7DLitWOqobMPTNTs1JAFA5JttmL4X+gyYoq+m4CV+hID6m3qvO0rQ79TSmiWZbI
0HP2QltXdbyXmrrP2sYorrd7TK999j6skDrZM8qIZqajRhgQKcHZn599npsjLFrP
9BkLaW26Hea2m2Yddt+5h0/nGBZjixfi1tqkVR7FOYeG8URchqNWLONg3cpZN0SR
Wa1qnyS5MdBMZ1rJz51QTQjmXTpbvdiBeIhNzoddtIGXOYY8FzfflDenegc3bpCF
zd7wstevFrgTeJfgm5ljWfAEicw06QEf6TNhfFMArnowjpst+yMJvboz8MBXXoGv
UM+s+tiJKPqTkXQnHRriVKJkenoR+rA3K+pFQJiIwd7BM7auujm3Xsv9rMUFvTRo
gl/AX/C4jDzOflSSNEsVRb6w1sqwNOkMiloeEds5/OH5zkPpYOrayQnBS7feNz6X
NOZ4RGxNjahhatFvbIJvCwUk/1WiOpzrmvUVBiIN+xp1mrQB0SBi/tMx4heXsRC1
9Q09nLc4nSo8qeGfH7fTBFSNCMgSBkTkbtOUxTrhdwHk8pd69YgSa1s9NOJChs/p
2HgpqBHxtjnNNOasPgAcN012NWySzQbGKdiFBjus43v3o70GBICiKkxxYmdgexcL
RCIVezZ2FpFkR2K7KqWA95FP87UVzt/bGGDHPVF3t4rtdZFYp97K2MZdX1I6tZSk
r2D2eZ63HOLBZxiCIAnGcgwJ6bC9RQnMfQJD/Z2rIsgUOt4xexeWlButKhuNsEav
L7rv8u1KFjgxIfAxtN66t3pEYifIAzgSu2d3xPIw6yA6GdsHkUYaDK6ItpLGzcB4
yWNAgowUbJ4BjkMdThHP9S4y/vJ3B+JSe9//EBF81F9gMCPLO3k4sfBzFgK9cJk/
ZPuj0FwKlD9lUKMrI6vkSDe4feQyCIJ0kYFIxiFz255saS2ZMHcSBhzr9pjbYWH6
THiW7ABFoQRM7me9r52+nHRw03StR9vefMDOoXIYEjXAXlkTVgbCKKgHQMHpEOA4
qbm48yzp5siH56wINFVDdqaluo+LES/eQVDQH/UgdhLPUAQpe5SuWbea5fHPgR2z
+KAeE7czyrQBjlqEGzACqEgsz+1bFvBO4Wfj7A1V2EjxSKQXkeSAGyPUcB8baxPb
5BFJgGEg4BlhQM/VT1T1e/p3x5AlwK56nTtYZQ9TiCcF7A47iZKeaVzJaSMWNBB9
XvFtgKZXxEhnBPqQbRZvnZvt208Zx9uZ+IKveHvm3G8RugCHr/hYjB60fBNe1HAM
oQl2ryvqM4dgjPo0bD7yMp7cQDiQ2OyYHDAYOadvmxyOKbuvldR68phZNSsIeyE0
oqo2V7UxFQyddIwht3MmqW+5aYDtZPxS8hEJLGCVXeq/ndow5N3kTDqva2Vr0iOe
sAxxpNT9vDQcWpORvkAIVeBOfF6bTJOlleiv3odk7oP2nfAkasQqtdr15XV9DLX2
Z2A3UsZm/ZNSoEAKVz0vpaPtA8tLn18qosDTh4q8SxVttYqb89iSshBUou2bF676
WXmtCQmwUPKErahOGmYJdqnp3D5Nh9OGGLlWoYUISW6yt+zkmq5Na9mNVXbh3s0O
YX6nRBrqw6iUuL/7smqSQl992vGjQbl0aAmG7jAUkKTMI9gbAc5YssDdwyRCOBwj
Zujjs/ktQbUvlTrxhGGsCKa4NW57VFkp8QZMBkLehjcDeeVmPYlHvYKiMgQzUXiR
iNw8Ylu7j9ADKPug7jHNSNtJPV+L4/C56Z7faaoI4zyQny3A+HEE5Du/Hv4WmpAF
gxmP330mJgC8F8sfOTBciLRTgED6e+gRvtq3LtiQL9BePYqZkuMBzLcVHa1+1CZl
3Hl/VRgTY9J2O/F0DD6ysyQITamHmUqawXvSPneCBgVxkaFJsqsEnvclQL2SjgxQ
rzcZvU988iLjQPA4zlvpz5RlCjDCs0eto4L21HsmYGiOZHCy63O24eWRmEP9cUJ6
ENfQvMXHaoMK3Z43t7g1yGP8uIcOCzqORfBH2RM3pQpstw2UfDEqAhbnxraK786r
XuTZyLGhqq7wu33YXlR4oG+WsStSwo7YCAX0HRZeqKdu6DXpt4GT3ssAB4K7MQRf
i30GKbHsVLxrV4IxcOE4uvfZvKoNAqzHFjkCc1ZRytSPA+5qXT01pbd8+5/8+Bxi
aEz4L0ECGno7VRJWMDViidrbHBhL+SHKPjuJJtI2A66ptN5gD+9jsqmK7dYxi80c
th2OpPd226YxBo6XSlB5WagKJeWmPF4LoJIf3czpd8QSxUX0L7tMXOARUJVZI9xo
U3l6kS5lgkYWHKtqexRkDANS8U3nCyPgGxf/VMUcHHXZOnXnhsB0JfDoUSTG+hvx
VV5sRv6bYbe8Pay86fs4eNP6Gd9cm+j1ODXiHGKzw2h7sKbNw8hZlYdFFjKLtrGo
OwXl+jy+bLKREAsrJL7yL/FvkKQ9c7xEaIK7+xmNFJ2slpJOpElt58ElqQI+9bn9
vI6//rIU7b3QvHDO0Lmjh5QUbMh5yo4F3vzjxKGTTZVS6qnR7x6lVsVhZtSeuHmQ
Jj5a1d2OWr+TShUrtWGo9/UgIxgeX1rTHJxhLMrv8B28POnKeqWrI+1ypHQwk1E5
RXGFCvbk02EeMstmV0vZTasrISh8J3D1RBpQ3deReV4nNSTY15ES1YPPC7zmvYY8
dTKCWcdvGer2dBvlpmSiVuLYhSOkJLB4kbaLcBik1nG2nlpAQhgB0S2S8yPFFLa7
eI+XJSVYNYg2Ayqf3EQ0Q2Jz7E+YS75PEfW3E41vdjiaxm7LwBtj4nyoIJImCFpI
h+FEyYCZIQhWw8PzV0Nhzfig/vuAQBE/JOiYexQD0fD8eWx2BnO6DQD5Q4qDv2p2
S8RxB0RbCBz5ihFXyPIyENt5OAnphji0Kcsiav8fX+he0sZkcQGUMD0dkOg94S3b
PWk5PLnsc14yNZMX/iTMGL5RAavEgb2wdrwrEnpenuuTbX1itcu7Az6OcH6/1H+T
ZTiNBT4/7eD6GMmEP0wxm3iC/PIC/63992WYveb7yintg0LMK0hL9RONQiiUXf9Z
sql9fgg6AElIomWdPX2DNdJmo7rCsKs8I17yqsh7MD+buIM6/mu+FfXXzWpdp33r
V6UNbDD1zbjI436rrRTdOAHfi8wO92F+kLLAHTWC59z46I/j6NYT42SojwwGqE4R
BEV6yLVH0WBW3eK6cXf6Y2RHydEnBvZwlFx1ChOxifAtVuBvn3ZN5d9rytz7suD1
/HTXGUuUrwsNBFeyMTROoz4LltW+CV9fdf9ucR7rnGNfOpBS/0NWgqEMUxCfUy2I
CJmF3D4ggy8oy27+BKTkJqYX4zH/bIOIdju63Xtb0QW8sqpXtrLyHePyQcMxtfTh
fDr0uGbJNx8KZyGojMLwLNQMJ3XyhfyqMV+aHLcPnH69CbC0LKDwTTgshmu2kFj1
E8/i7qGVQ0Lhny0kbTkGlu0v2lRpCChYqJIF1ksRk7G2dX/MVZFNInu24aXvKHtD
K4gXLtTxF7E6SzO0pXA5u9SSaZr/iOyEyPBKBfeKiYcmmZ3SlOwt2RRftV2euz2F
I/RjU6Hfrzo4ZAG80Cixe0FyC9LFaKCbsOlycC05qNltiQEidAW9nPnFhVFdk1h2
BqN/J/eV6iMuxi5BdmhBCsVm4h9hk1iZ3Dhuc/yrsdaO/s7YlLF2zez6PjDybwyd
fWfjdFCto3oh/A+8s8YcmtI/IMJt8vWvye7Wk9qwZtsH3OVz1oaxtNSnBeb7QvZC
HW1kAKJG186f+27S9McitCTDxcYHnBhTOW/ERWmt3aEGfY9+1/bFZINKrzfXZFjB
6CHA7wACzXrfzptYvUCaZYzaDIjMS6Bh7Y7XeDus90B4lAGXwX9GH0M7h2CMcH/a
ZgKlX5A+u5RUV7WeA8fx2s2kngtie28OEnaPn4hqWIi+mHcKRDNBpNF8DzPg7F9P
iGM/tfyeuf78iaAwcSN4xxVAZiuuB1+f2+h2kXDebGYZeERjgRLrKngKVRd/dgFK
bgKl08firmxK9YCdSJF7D49vykNUIvlnIEadiYgxXJDQk9P9hDZNY0Y3zoQ5CMp5
PJFguEA732c7BiaCf2tBasunn4mgYSdYP4jl5YVAp567K2TS1RhV5SsVkfpzfsnC
bMkSzOgEgG0cQ7Ulh2kq0IQ1XB/lfSnIFWk2PKu2qQmt9GxepLVSN+9a1FPg8D1d
yJZHiaLDX1DkE/zA4evi8Ll0RXXe4LMusw3GcL+897TinpvOSk2/6mby3O53a/p6
odN0BAvRW3JOi2spUydwf1/pjfqjlNXTd6zRFEqhceik7FRK5oHwjU3HhyxNZW2V
FNzNExOpDzGTHTat4Pw2gzn3p44S0FvLBegulf9J1kjYqBxPVWxqk14MXw7acjoi
nOjHtcZmqVijzQqRFmlJnRr5PBEzwuxRGaYRhFM42po78r+HsO20qYATQ/aQ47ox
PM840uyleHkQZBcInzWuDPw5EbmBb+yK5WgIgdONQxbmAaF3UTenDdwWbnts2D71
DJQsLu3/HNlHmxFI2j8Mk6RI87k/2xOc8M4q4OA2LaUGeQMLVNUYfEPfRqhbrzS5
WqsdJcMVU29JEmqJMtJn74Cu9yDAWnIFQgiWmVLIMyVz8nnTKQ33SCKuJhefOYE+
Q5EopwxNtf/EPnGuwizWTTRjsJ4r55BUNSALnOvB4Y9AqaceW3ZOcQcp9GW/zVut
NdGXE+VvFSGIcoJ6Tstj7zzjJGTJIOks1DN0d4nOsUhmVL3nNZ2fJCCsZAepmDy8
Dw4vL3Xp5NZBwj0FasCSWTUvibfszwz7tljaSznLpuecH2GDU00702AhcO6ZR1yP
HUam/5sjm/1UtRG20RJdOMQ8vZOrx7n6Nba6IBgg6PDyAUfb6rSaGazfx9fpR7c1
t0PmcT6i4q9Z3hWL9WKlL5fzu83uPNJlbGoumfoyShvOc0K4dvOUj3x0XBA8nJnN
nqIRBkTDanJ5j6AeCK0ioj98ETsOcIizl5Dumcq8e/coqr2ZMqh9Jj/97AToxxlw
oJiIKAIjigfyr2d0MBOVvHLJoqOGmmZVcTmQJGghPc25daOfzbV3AJYmpxFq6bxZ
r96VF7ahUaqS8iqwyE6bgDcPoqAkKG5kSr3VozIN8BQ12tlRQQNJ3BiovIA+0X4l
/v74ybS5q2hsrPoC2hoOSPZAyt+F1Rx99jwK+W0e0Xqj5zdEktIqfQBBvWQVx8rk
UNF5qFwZRf/iuMsJNjZMARTX1OYIUh0fFu7NJjHpE3GcbqkvCN9uX7hGHpQwYO/D
aGuD6o3IHcjUj1flEQr/0kSE0A2bHZGhrGXqe/8pL3W37kpSGkJnKj3+H66Sx8rY
jC9lZW3MXlkRJ+d1GbEVaS3JD6T7u7Ve8cDczgNJWWMJffXuAgIj6CCN5k8wyQZR
4/C1URO/hSv/GEy0MkyyxA9LNJ/gHLkSopUWoRoAi51AgL4x62/TvejUjOLUoS5T
6zkyhqGcc9SL68/sX33jqFv3LcE34H5FK3fQb7b91qdTWFFrRJE4k395IMvLNdQQ
m5yrr3BosWFC0ZsbOFIE83DQYZ6ijlvRBhJZZV/4PVSs/Xz1xfJcbNYwyY6hDHdW
dW6umbwluMpP+Zhv2kZ7fiKRPcqo2TEY+MwV1ZjO5PpEbxffVALw+OFEmnbe08B+
F1YdHGzOlSSRfGSKehFbry4wB/4JAedOEm5MlKj4SsSPYaLGl1rMP/O2ZqGdIEgq
TaLoRvFfYLjiA4Dbow6hthq5Cr496j7sFp5pxq1CD5ec+6MhRjzYlSbYnSdNBTeS
ZV8+vsmeZAgr4azfTLUAC7XNCsb4O+VCm6X72+Twa4roP/v/qf3pHcla58UGZR4Z
r2ulNeXVnlbKqLwmbLA6InXKnrB5rNt9AWcLl7tHgzAipyZ4sn78lgvil5fSlDG6
g/+CvuvBiGzuUqiywqfF3r8o5hc72xiIAn5ZR3w3yR3ZvsEpQ4jrOoQB/hELoCMD
idxNQiShVKfsUtLSKapOUY1m7X9BXB3I7Ht+Y0638HbWi7E8w9dTgeBelONr7jU/
q4EsK5CpEm9bCTRevNSDpPRypdauBX0aj5kEdORev8C+A3AFlEkdp5HsuodywM3t
gvyXtRBFOZvdfKIDgEA4h5nFRX1i5cFyM6TQB7VBnIwWcLNZ/C7pTNpVnRhiJCHl
takdLfnnUtTHl2OzEV4qGOc2v8e4G180wft4nwO/iANdNT7OkOkE4bO3vBuoEhsY
k4w5ZjDD6DxvK992ZaTzGXq1HlsZ1HMRuJAVLLWeF7uSgT1WfGIJMXVnDtt8ZKVM
iEwY3ijDY3x/m/0kvvPhrpx1iN1M5P188rmg1mAfjorEHG/L5GiJm6U/F/S82t+q
aJ9lANUhVl1vyn+w/Vj6YkkBbegc8Ij3s1AR1bUYqyMYdSII6oYUmjEvrQoGlwnD
8/k6NF4kOeSRzG1OaxgbrUpVsce9yzbesIRnhSRHfXfz3PHOgeqcumMNW12hYlOw
MAr3affNLSlynk+UgtFEhQ5lwu9KSCqiuhyTOmoBoL98wjLQMuPjsKxvbMykW2kl
rzn/uuvWCJNCFrDEGz8/MQSWGGMl/xGntiXGhEtntHMz39CNc62UcvZwTCtUWtQM
t3sn/hb+M2JfLSBgUTHCNb4cApFy2Nq08Jviu9Ny/zBQNMlwEghzr5TwBNQfRctI
OwiFJO+dY+CQ77zTIRFs4G9Xg4dkIXmzWnzH6BsD+HbghLQUVv3sSqMJBi8bblcS
vAFgKZfw4tj8gEcYo1v5vRxTfAOhOBGepAhgJBSnOUbvF2Dxl5ZwpKkZWbc9xsYh
Felx16JE70N627fqeuScws/BdRMmQf2uWpZUeJFXLxBc2NqHcQ1k7uB6djrNs5d6
yoVn84FxDD89Yy3EVow8YUC5LZUkiKFdMhC6yDPjTBf02aZKlD33WfeAPw/9StqL
/VH1iC75Vy+H2/cIiTeaSgOU6tocjkUZh6NY9s5ZKetqYSiP4tr8B3RERbT/U0gp
dLD11rTf6KnqeuysLDioBXyxxTrYYnQzF1qkeKJj3WSKQdCYfkTbkRaJM2/137Xi
LC0wddPGpAmruCqh0eKKQYCN41BrR7BE3nRP4vxI4ryOQsnSq8dNmjoKphyg/7JA
7shETLmQZPmk2c0SA/O4nJERNqRMAOy3UinnA85U0tp1waOTVJq0OCqrAxLQVVa7
XDWN1ADpnuS7vuoTz24NacR/q113mWZped3XIi3XU99AReAgMK2GVWOXhTe43NCm
gbYLCp7qG3dBGrMsLkbfe3gG3LmRBvsfdVqF8rz0nSvoYk+GrK4d9EU3iY4YWhw6
yza48drLqCW+vDgDeB8LSNA7YokUCX9l6wKzJWn5nnenZuDeLUlo4WkSQLehu5U5
4Rcxu8ZEJRwSbbpc0gJlD+63sEyaEIU8hkIx1H2JOrBAy8psolA/djcXXDVw1gGT
aIBxqQ7tBN0IFr5ih5xH2ESGjaELJmlf3918QSPlOZpD0ouQRb+eRa9xx+8CAFh+
uxvsXRBEqRBtzJ/hRH3yN0UtWDKjRRCx5cXhy9BUGF0avIdry7u2NL43LHhKYnd3
sUAgvfTXulV8o3ymLJQAyYJVCimTCphokaKlJNH1ncoWDDV+JRpyE9H5/9Kmvlo/
uk8CDCeg305pSkiMLmYftZxskQy6jA0WXOZ3kJGBxSeSUf9787uE1WilwBlsWPCV
nH6lLNqGiNGYy+caoEdtO/F9FRgyjvxsP+ROjtJVs6xzpx0brGu0TXmLF0m66LPD
1pSfxPe1OEW584zDHt6CEdKm8iWE7wIhp+50gQs0c5i3bw3XcCO1xN5ho1Dsm7pb
aKUURkh2m8BHVktPsxtoJ2fKlgvkh+JuSBM7oJ7mBB76PVqheHZxQr5FHwh9rElp
G8IYoRzXSRk4PyLrMt5M7Z6wVWHwLM+mXEO3ki9xmrtbxUiTwGoE37dZsQzPllzx
8C5DN0ipuLy8TNGEfjhzActLF/aq1/Gp+LxuDpTv+UkUJ13EatyzfwxkX0rdxlue
YrrBDNCQrvNtn8YrJfS9RmCN0S7cmNA/vF+tupfvQlIojSwVvt/FaXpRFe6nGafK
r1RbXAqykhOr/2cf44QXPDu3ba8jb2Jj0u22TmhvXlQqDCRrBmBcqvnFvrhUruSU
Ii0SaD2/OUkJ9T1W//48w1aLI/hVhYX3Xu9a5vb+g3Nh/Dp7t/oUJJMlldeL6NRn
AXQJMDmuZ6VzbKNQHIqNPvEU1jNz1cGnjLJLr03T7nbV2eLOUPl7GORIA0tnPL8/
ALfPQtMOHBDlaGPWK/ZayFc+PTQhJz6i95ybvAP7em2sQYyQbmxtQLH/DgD9azn6
8Zvhan0ggTxL/vFKyt07PyaoBgcTVWfstJdW5NHK2Fkfd0+VeOxFCQg2NXiFCUVz
LaIgxw9rdYpHbdPYy9xOY53RVpuOcBPOcy/fOIPOEiMQt57Ept27/1+4G7gKjrTh
s6KPywJlboTRtgumvVf7xBilQ2egZpkZ9fT20KTKfnvZ3dMQ5uDUn2m/LeKkjT4l
GLMj4KiowN0LiDtTf/GDSMBvQ/cMGmcSkJkcbkoeRZsG/Llr/56LWwFAjwLzAnl0
QzOPDUPiKzJP/DH26GkvRU734N4YoIaxV7uAmjRu8caFt72hc9aSbMvEPeW7RM2/
ERpIqjQ0YQRWTLpj3IxNYBOptjY6/fLO+a9kl4BiP/M8BS/56M5Rifz8T+olWCXq
8nqZ84mlcYbalkfJIDuUEbXfqHR8YFXOMooQMsi7RmWteYUg2xsLM+oZafEqni5a
S0q5AtkUejiH4HL3lRbv5pDvclNYBmYkCMpRQwaz20Qn1vrLOlFq4xXcZqO1DMj6
2JO+CqbDJgDFWojw4udTr9YtpyqNY7q4Y4BBIq18tT0zmOCzWtV15n5hyfmswnvD
N+/sqWVHuXFZMpXiy8IGHdPxZkyxkyeyNwQletUzAm16QCHI8Tk+MtYdw73cN9M7
dosGh7/ItduyXex1DLw1SEJgjCM0XYwrH0WZEjLss8/hFb01yI72Y37itafQ17dD
mEhSjSFIg5TUQ9MMNXeO+J5+Z5qr0s5FuVKsML6fNr/qukNiWjt73L830C+8OYq/
Dsd9vTmlb+NTovHrs0stsx+iqphXJXO/SKdv1on0IdRznLmdzqnBlWDM2//aXpD1
zPpRTIlQay2GycscibjaoPaoteKHPBfkR1DtGRO7Yy+Fs58qyaLPDWnhEkngonzw
jJxKf4p49fWxeTE488/tyBOo4h9fz+ZzZ6mTahSLh17/1pTrjDLAaE+g4eIi1R6B
iRzrYJe4B4WiWFncQLZtg7L+IsxseTRQvK4kAoo29+g0peyKvwruCVw3uudQ3XLv
w1wr4u1en+0ZSd/QR8UBQmu2Mi0L6Q4FSdW+UUPgb7I5A73Wj57i5dyekS/G+MBb
MBb3PQkT9XPsfjWXddbHQJbAD228/bQX5yV26wGBAPtNtd98f7SCD6J9lTVHS7eo
253s5eTcxMVw0ChbkAtImfWUUjevHtbgdBJNHuofNsyzPq03dekZKKKKovT/1awG
hrCwAWUN/rjmt189iJjvvyu+eE/8YC/Qv3RyXxw5+lyf2p2zW+T7n4keY12YQ/8s
o7h/qmoaLWuK3df0O4wITELtMpmFGWOPyNGGMy6raHM7EN4lq6P8q1bnsyPqOmsh
tPz7MjuW6hfjC/+Iqjv35HQyh88b8m+/cu1r/4kI7+d5vbOwvQzGHH0NEnHc08W0
iVY+KUR4EE3KM8eJbIX3tUGLSceY2DrBY4S1+1MEY9864Le/HWMKoeZhshHjW0hz
Htr8OcqIYVjQlY8CC/isZT/X0e1wK4viAw5gcrHt+lETP12AcEkowK6M/JaOKF8P
1J5EuQt5xfVKt8SzbfXHQ+IB2gfhWaiBkJYUrCOf0qCfAh2kGXfiEtOZJjpjZqQB
wH1fMyGUqtnqx5iQT4DRamAOGf2ULNLt4NfiW61x8XabcZaXeAG9zmoWXD9U6EHZ
Fii5rYjwG5oAZ7Gybjt3Tz3u/UAaTyTeRAJkaaCRyOWx3ysXPUGE0kxTP3N2NWGT
0LWrDO7rEZyhGByAEiqLsD59E002WeQdPuMEDfAbHtEVP7aL//z7frcNlyM54kxs
5Ttq1QdxMKGfBDDT63JShcanNmuYP/8cw6GeDbbeRp6qb8OH2k5DcPJWaQzKW/dj
6nJE1DhWDLxz/Z175AwrsyICmaDz77AUll7VzhWLkAdkxgmQBgkW39dGS96w9KAm
sAwO88WOMkpKFUnX1eM8ORxcOAW3/XQd89juH2Wp4rRYo+PQ1iKizZtqDbR2RSvx
eSsZ8oOqgrsE6ZKy3VmTdIb7V8OOlZM9K1eVTI2APzVOf4WYVZNz6hmxp3Ug253K
J9FIHDhoVSeb8dy0+oHR0Z1vIgLFMen6CpYvLVDJhB6HWTRdgeK7+10Oq+t22uuX
QPSZqX/kNo125QdQZkyDCTYEsfcCJLI0adVMwnR5deKp5WdURZetM1iCvE/jj61z
arN2Ie8WQLIUJf0Vh+JyjocXH2toeFhNcog8YPaDlhg3Avjef2ez+KArFiItJWls
Q6usVvRydl1YoGFt7utVofHO1Bf+ImMEgqbGpMztMbrlEx5bbmmkqXupzK0VLt+r
ZEe0IOUWV6El9OlkW6kBlMCyf2/TfSX7ZWA+39YFv5nyb5zn9/jS2RBryTx62s0c
ztV9XePqXIRBOU+W30EWcXDBVX+oOpvPxIwfLPTkaozIJbm21cpG1trGhTzbMIzs
WYvMpUXpAkyIDkbyLcbTS1n805Kx9/ejHwpPP25k13Hq1v4y0i93yFknoDd2PTgu
J3LctZYNiBA1JBKpc8MjLFXA7tJRiq8KqOzF/S9GPoKZGHo05tpuNjgeil4KHc8G
bRN4Bf1Lzjohma1e/uoYwLF66Dx3tPORDrWnQqVr/DzPWVLqZzfJ6uus4s73PlTn
M14OIjnT7J2OW335w+ddhy2/ok/5VTkrso3c3ZHRfFEOB5pG8QVGJDMFU9awP9ID
vxHQkKJSv/5BpLqaDIT4JR3ppBluzCz78TB76eeRbi8IfsDIQbxKD+EglL4qd6BX
NiKXqenLYtKw10sSw2zFNiR72Pav5//SsgpU56FfaQYSK3R5ZQstv2NNYJp+sYrN
HnO7JoSJPofpUm6I9TE58ZjpxETCixED6Ezx9A2q7BIccxP7dyj6pVaa0eHX52Gr
IGNNfx5pjPPcA5QgWjv6W06MPifmMWLvA+Swa+7eOazjHOwY4N7oVLjABi7wpVa/
H2QiayGuv0rd0pGneTtnhuXGkqRu1Xmmg9xIFSww0GwpyOc5ZduJf3ifYuiJ9hyd
/7mQWMpRPfOq2VhIxeSpG81SIUrZV5jLippI+0j+BpxnE6fvtJOHgzucMNo+tIoh
kOwGOt+jE2IowF99VqcxSAJmZq+AMLdNHjVKHBVWPZhyZSIve27WwvyHlYI1371d
fAK4P5hNB4zKi0N0tV7OYg/IKX4FVhL7vZ3Tjj2P+rasFuxv1KNmA/sE+PLCSWQF
v5rmXwhVAiRh31XEhi8zBci2qTRGGMKI7kK7aSdnwntho88SleY51CN9XvZW9MoP
MlFjiusE+vfx+kGsis2B1vzwGVuohq8ehaNqmGuLXAWChPLbKm2la0uQysEwWXB2
m8xHbxpgxpEM+LmAschuxqIfRl805HKLW+pJI+tU9mLmQD7LFR2Bpc02jACrNNN4
h8R0XZX7gqLzGF0s297B06CdiRHEm2LCkUjyau1jTDoNaTomEeCP4d3p/erU6uAQ
00NPXUORK1oA23fOdBO8nqfwgvqk4do/cehmF3Xv26Ee1JgY8M0UD4ApDRuHmrlp
86yo0ZOF8lxE8QFqJC9PCZ4u15MCAHh1YcPeQKH1jZi5lktw29ZHVT6LhT4lFvco
GEC8ctJZGYdPSKkd/KdOBPq3aKzuaRR0nRnHAJr+wt6Qbqk39+EYRJuMWOadOpYW
ahJdtpYxWMyQyZ23u9CFQ+dy9SSEy15I3SXBIUGRb+WLoIILBXNessVXK4jIPAXu
QWYNfggwvKEvpyq5d5rHL81hOz49bU3voeW/gb3o555wcjq8kaqX0KE0e0Zr67bJ
vN5/OeAn7mobd1FvZNJs+Xmu04ucNGk3j0PaKFAcss/pghiZJB2LkgKwhf1oCgKs
Hl2JrTRXg/HEN9dLPflrhTioq99W6wugkW9gJeZym9e9jiDP9QaI+C/4SmaCgBpU
5WfoKiKTfLWI68GyDuQuQjEWYZbRtDMyaDAnnI5Y5FYQVwr8UWCVuQ3Et6U0ipPZ
DdCPbR7GgfcHYDpn5on03ncI+uYsp6w3BXGYXvmR+uS+KiNRUhUTjlB/ZzUAzYbK
eHG2sBfuu5ef+5D4A81GnDIi/LaONfia+07xm26gpmhn0CFSOYoGFM12UGD3nAvx
EdQMx2SMNHfrGh/XFxTU/u6ua+46CaUOuTIO6WsKa1buBfjvKGU+W3JplLH3icOu
moKxlODEPjpcc9WoUTlVlhsIHKHn8z0OXLY66bkBCU39GMQPTrta8Wedcw4MMxyM
4BRoFcJH+bkG2eqQjIifU/1bvWi30Nb+Zb9mDCwVv+2rNZX91lEFrdcFPXmIr8G/
yZ7IoVMR8xOZZuPbOHlVQXmj+segmWksfCiwnjuneCiS/cn+XI2JRfMQlwjSr85I
FniERz7Zp8m1hE7M+nqwp9hOkAI2Wd3U1bE91GJNKScuPmKgBcJNNN7qVKzSts0B
fdZbfqc01uVtUTMHYdXe0w/kNulwIXlOSwicnrdzV1r2LeGwk0+4XSAjB1TwzMQ/
tuT9Q2JXPf/5ofvnQLwovlmfRR8EjC/BBjhEwhNJUlr+rFPP3p0bVK5OlxoNSkeL
hMgpn21+x6JP7GkS5BJR75GJpmqglI/EhqXPd3sD/idBMkKdYOtDtU7Qql5tSrVR
KoDfE2b6SC3RjdyPcCp1o4wbnA9sPV6oE5Mq+Ue0mDRMvYu1lkcS4BZg6rSCGYh9
v/aY3FWL3Z0b8ttuuqXCUH1IdION/kB4KIPTqxE/csK8TZ5fsjRdwyLbt61qwlLO
0HAkIooeyzV76VgnJPMpUmha9SakVmJGzN0AQNL+n+z0RCW+ghC8CWNwCHke5Gdg
If0cD1h65gMvdCedEdiMDrLFiaOGnG+AphgWIMm6kmmG7+h2qZf3rb7uNxzKyo/t
EREkKfvUzduDnR6QUasdNxaYr0HQ8tb27pEjtKRDHqX3rzF1/H/SciQcjlUvY/lv
YKilqIbS/OJS0U0f7bpwZ9nssSwEBk72Iy9kNJmuyB8olrOnqoRgAQ2bRK8ix5cB
GORtvLiuXSdye14qDtbH56wHO9x/ts/89U4U3v12iBRr31VhfBlbFw+ndfP3V+3A
miaNEtYQUZaotTaD5YsPJY++mbXv9R31VCTmq0AV9e3KTzgFyBhh8Us/xXc3+Q93
czM55x2kPVFM0aac9O/9AuWsA5S4ycZBEBA/KgHTqmCWKmJNpUUseIv/tfqPcJLu
w2qITtCvGc+A+yQc5COSl2w1DeDAp4vpYB1HOiGiGc4rJea4YDYtoa7lByimtiGN
dr2ZSSxuXKUDK+rqirG0jAz9tq1/wVgpsfLvPMZD3MxLIFgJ3vDMZvxWTRcvWmzt
SqPrgE4tx8t2C9zdeJ7gizZ0XowlQMyYNWPN1F4zNAK0IzbXnm6OBTPrrS9Fp7gv
XnprHsH5f8k9OIVMfy/f9pgzV0kwpeHOtlZvdTPqNuJcYQgdLJrLybh+EsmXTywk
PmugtJaFcoNERD7+VbzE2ADsZTqLPNwPV2yAfgLALjH6VmpxrWOkJunS2ytWPr3r
Dq1WUk2OSRFEcecl7d/LlZ8lftA7WB4KIS8OsY9LQOV9eMFhj/2kbn5AhSSRvsmu
LWpo5oJ2iwIHcPCcaHFz1vsezRBwq123+l4XvE8zXzEQwf4GV0WdzSBkNwLHUy4k
grBSjz1xGKAx5Nz02FwoEOXjQXjk6QrtX6C3ch7hcOEt/nazUV0UxLzbx9JgDVhE
uNfEJZMuz9H/EvckdX2rhP0Hbgdaig1fFhsDqb5/YUSbTH2UFjehZkx5hCFopkBJ
td6oLA2/WBbBuGTrzigFmPFiIx6uZWusO32xwdmq9aHZRaRlkaq4L+0v3ENdZhzt
B60Eb5avBfAj6zXQ4h8FDMPh0Mrfz9g+aQvFlneQxU6sJNY4ZfZza1MDM6Wqh5n1
pJkxhA6Fs0BDfdAUYd0R8g7obHMRQ7CjZDieuQvUczV5v/NAjoDD6mjCKQEretuC
ndda/72kMjuq9gMrZ878TNGsq/3z8Vg0cDX+TZqRqcjYz6gRLWc67JIak4wUaFOg
MK2p64MgmncTZbaPR/snFpaojfaW6LKVVlF6ToOufFU0bnZY/s1Q1zeKFeOa/1sr
m1HHNH+ia7Y+5sCO2D5j7dkf18HHoLsGVeiM3PbNwc4pdLqSUErj5QoI5DaX7v6h
prgHUB50KqLpgo4Z+AFyfXpntd5viQBFI8+H/9LxbyjsOtXmCjNlp6151jjLyHGi
KwyX39tK8Zr9C2oyzXPFUHDtFIEEA7eqkR4UFCKLw0Oyk1FSjdTV4USgWGLL9lNz
z+N8CIAXm1P3hz3X7flYrP4lSgolkwDc6cRo59sv3dsJi/aaDnUKRTRJ06HhGSy4
RVSza5tvjWLZ7K8jxKg8FuOsPSL8X19FVfGz6OTPATCYsuY60aQgwlY3Uh7LTxEs
rshHuAV+Ty8I6WOfqe2A0Eo+9tScfOtyykk79wIlnjo3Nv8eARnlztAsNqZUl7NK
INyjW72YWiGAu9gXgeHmd54/maz3d1vPGFexqFGmPTv/WyOmYF5BEs+MpRvvKMc0
OkY3slcbPVAR/O6wJKVy+j8tVrGMN3L8oNefdjP0K/VSBztPo//mM4U6je/qrTnf
lIggaIZ8LntJdvFgBjEz+cayF7C1jxiXi10Pfs5n5C37Xkol42v8dGnEeYE8yUmD
B+VomhFk8JQIc7YPPe5OpjQo620w7tG1H0lXP3xRZKuxvb6qyWBA5nNofriX4ifq
Z6p/olboJLN4S23Bhvy7h5q2BKM6KYXatfyf1CdqzJZOwQcTosIF6XZ+uy3FmNxf
JLVw7I/Py4/nWbqjSgqyOMF9dn7vp2CZm+JVYe2eHowhWmJU0u1NWbblhvTdzXiJ
/Z2mv6Iy5qanKWYSMXFTVVk7VMe8oTY06uaCTLljQcDXLXflYiHlbhGgVMIUapC1
TSLuwHeEiKDepSkH9CGzeYEItIv9FlH4XV51lypR8picmLldflaUfK2KBT631Qk2
XAiJ2kP+0QUfVIKzTM3u95JK6kbxiRa7OMNs2/b73e7nG5ddzypJccbICZBbiNDA
MzzXJwrE24nFN41NJ+Ajy/F3AG8ynH+pW7sorw1MJp7e4NT5G3dnu8a2ffHfTd1Y
+pNkzCgt03xAzZ8KRHBgWYCEkGLzhFW8uiTqrPUoQ55e23GPlW+2Ed/y+57+q6nx
9eVYKL0vXPIGyfrKAO24PBVLmg1+UdtrJtAchV5fgMpLDWr5PKfHyJvD6Q5OTGn8
Ts451euOIy9toYNWdTACt4Q9PBn4MlTbxZH/syFqCY78oMubH7oRx9fIgccI1Pqd
SaZhx/gLWzWZ6qpZZx1oKEIYHmT6z2BWM+/vizun2/iUgi0dAwETSASBoHxkrWDs
6JleElcSAAevlRkf1HpQFf3mkjm4yuo2nXu1yOAfWPun/BZFb57moJ6z8DVPF7Ma
TiN4nHqjcRmGgJt19g1QbTzYm0Eb6y4AGnmCOMdr5C3EEI+wcH+lN/QAuYt8QBvV
zyxdVnE5GAEyoUB8GH47uudNFLOZf6iu9nVDa/8inhl5KZsxyG6ZCiF7ci0CfP2J
naKq7hFfKowwbWQE+8PvjsCpYOJM30I5JmTgSVHKyKacbiDffTcztekjyqepbcTo
ukl3QWx/iCi7kx7hsozzfh6uH92MR5P36pM0D+08hTzgFqGFdCp1RUGwLgVKs3wH
/lyf7+0Q3nsti2LNmM5a6xi/7SyZdYIYYd/rSNNo9aSYFZ3XvQ57T7amcWFdW4mD
MYdOFniaya2SP7vL3MKOnxAYrdtFVx8h7hVCWvDdElQett9sCDyysNyBX1m1F0eY
9MSico82aVROhj/3Cbk7OzKPpINx2K2Ov+sCCxZKTZVoH2dxoIHDQ01LrTVMRG3i
u0utVwTV8fNPP1ry5vemZzcTnCjDXeV3R+VbOq0ifNeedBMnTE9e5f3bBLV37m1O
Q4Pf8ltNYxLy7iNhCMt6i3kemoBbpb37v5U5Vh1xQ70Q5UDir+pt9r0nBoQuDOBV
by8voAPUZpgufqj/Js/qh+IfymvAyjykX+4xboWmQm/bRzdZx5X9k4he3nCXxymM
ypcVuftX+kM21hvC51vWCib/Arnz7lrPe6uddCXZ1/hTzF55ubpxOhD4HS4y5XM8
Sar3WcEdVx7gt8yBy9o2M46SurX6NXWwn7+9NnVFgo5iCKU1izT6sShv9p1umI7j
I8H5ngwkzyn2Tv6qd+/SJ5a4MsdLItE2WqU4Rqq7c7qbrBigdn1swlJRsLFc1Oht
VLhryYOp6HRWP9LIEh4h/VoOp8PSC0gR3DsInf2r+jOjnXvZMFj1fDsGNNOQhpbn
uCQ4YD0ucHCCvCtlyn4WDKpGQkN+Y6IieXZc5ievH1tAoGE8FQd5VVoIzzXCj3WM
/gS2yCMp3BCUFNN4QrPQc8BHw7mN0HFRVRZoV21ykzHhiPhhVZ6WeUrZfg0BjEtQ
pIJzNKAwDiSVlo/N8N1miFV0eC/xR9Oo4e9uqI8NFYdtglm2CoorNgudOrRBdQND
hD/Vf8e3N0mJazpl8WCF+4dSJIM2mNm0bV1i0ZZKiZaQS1GEWhgwGX630RnS6aVf
vh/VJO99LJB/avhyJIKuq31kzMP87KtYxpO3gIvuMdjMrzDjBeD60THU95z8ovE2
Y+Hc8e5UKAiXyqOreJkuztjaAS9LJK3eKLi5L3K17+ZqGhr8Yxhnp1eFMzOQSATG
uvhw7KzbhhJ406+W0dLOhryNl/9voINETshOlSbUeCyJ9xwyZ07oX7bkN1AbZM8W
D6fQZi3mW2ULwnNkNbIzGatJagAerordsDnyiMRoFKArRL/+Wa0A01CTYYXYM/Yo
2mpgf5D2GM97y8q9VOhZS9hoXL/2Pyy85g62naMlvVB+/m6w/Js/2w/b1UABJUbq
4JtWvOxmLYm8SVjhcj3BQf0q4wbBLONIooJUVXDAkU3o59qgvUUU+WWJRovzhDek
H++F/mqULFN3p4yUPnm4Pk66AW5/cgVYRzal6cLY0qQyU98GebIirufvg+hx6gxK
mYPGncOU/2ybsMcDrPACH5aDm6dTRSekYYIsZ5K/zfxgEsbEa8M7txGuGpaOBH9E
VLz6Trag5l1lYH644XmVJKehbWzw5Hb6V0ER+TNFzXsrPn1PFRKx9Yt+AziOayrf
O/je/TrgPu5dP3M1m8rdR/5gglBnwndqLvAZabG2FatbolMQ4JeShSxwEcmxP+zv
pp63yaidio6ZGXnkbt4qF0mHuQqMBoaXF7M8vWvKCNN8B6JkKoVb3/paqhFqikt4
OzZ6YIE2FFfgiE4EJHFGXG/goW+3zP5Sx11iREtpX+9fcLl4jALXKDV8Q4oOJoiw
zFRi5Y5huB4Fsoz0w8Zp6ft1+3i2nzsKgRyewn8xCDwZsqypPtFTBj+MlnW5LdS7
u2J5NCr7FzMveqSBX7aLOwEpJBbwZ37iDE9uA718M4Mt7aV3aAee3/kxGbUiUZUz
cAxlopfJncMDlk0p0foasHvgtYbcieA/caXesw42FChVXksgbm2EMCHMZEoQaN3F
EjWLhjYjnG17gpWtE3ck1D/4BS9oryh0FDxirjkUs1/duilG5ucpVWGUXVtZJrzN
n0414ikVKLG+b9KmwYTrsmbhEgPKa8F+m/PWs8srsqaFvPB0vfzFzFasQVPBCyJm
G/bXKt3llrhAWSxVWyZ6qW16EYqCxQhKOMG6VmPfxKJT9N2Zp2+Y85zpwxgnOdOy
9HbGPK15ZZRaIAtgcxHzDjvJE+LVfVBbGFiNBfC/pEyc8/ork165SXiyjwp8V4KG
slZPi/rl/YhGF5uJ1iZhSg00ttyWDm9tsHpRwIr0FZ5UxNbGNBefwfp7WTPcsGsQ
vTgAkjDqXMDocpsbIsdrhuEVyXmy/pAPEY7q/LWujeyUnEP+6N+5aRElpCC2G6Cv
sPjYxkBG0kvhrteiebNp52n9rrdfFwbR9gOV6B/6vQUXVEaJi4VOFDlgWcHuEf6/
EGEpy1/aLC+suGJsgVAq8vXKrkioiG3CIK+4chPqoGggKH6ihfYh2t+oh0QMCsjl
txF7Uqv3Dga8ih/IhHC8Lxlot7+erUpgnIhtOWkTXUXeXA/urG9Jpxtlc91Nh9mP
Ub6EyWnRlCYbtRWE+oiIq7Q8Jd8E/4HGGrXJ4WyweAHXjbVmVvun2GcONXXEAzTZ
XNI+8ZfYj5eIN8xERXw5jKMisrTBRiUOurBRRYxMvLhWwOhfm8n3lvNJ1faATIAQ
wTsE4Z3nKyHoogx4z/I+VmOWFnFb/qIufN9rSbapWKyK7kd4JIKEZQJfXH55xpZu
OaQmMT3niqnVbhEaVBl0RQ/qDkIx7bHmjZRMxoxG88/rMfAemfOqqYJ61EvwaZgH
yYXnTy42IIzT3har5zPn2UADwWol7mtFhm1a+M1ZJ57DiIzc7IyMfze54AzynZ3M
+JE7xAO2453v2S3z2d5OPdoDFTycFQ/pn7wRHINb7WDQNA38H+DWwYla5ABJv/xY
XQcf3iEvJKkoZjY/AbEU6XOvOGvl42S+3LxsgWyT+5vJOglW+taHoIWFcNys0dHA
U9S5tPfk67c5tnhZlGcvo55SWW1KSEBQGpz4utITiwfLIgHjGwQ7SS4UTZNX8Kpk
7t1lxtXskhDirDka6sM9URVb4cAggSU+zCH2OtOoX9bJVljtt3Rx+CbiC2FpGsXA
imAgEeFncO0IqNPMbpC2TLs+u40q4Y4mvCMkA27kHMe64772RCHW6zybrqfIFAfI
Cf143Ui7MWEMPr1hI8EZFDz2VG/MlmmbP5bOpG51V4E43Zc573sZp//wJmS7qMP2
qPg3JwzG4hzuFqVg0WrqGc9kwjQCub4xmSXZnfbKCgdIfjbgwz4JWMok1iQ+LNqT
QGBSmr2KIkOWvX2nzMLExa5zKECv/KfhU6hTHOOCCemNYVehQDUL2BL8Cq1fU14S
qbPqtE5fhsmlc70R8X+daydp5QtmbmikfRmm+sMxhxwKDRhPq8zwDZt5N2mI2ooz
sJ5FBnMMg7lfgZqynnK8Mto7qpm6olyxG2zfM9l/rl3V8fsKKjfZSVnl2n0oEMxJ
X/Z/Yxu/lP3QoEolqjfc0yVvQOuqNlsJ0r9aPSx7hCrlT/KQt1Wuy3anaQtAhEF+
OEArlRaF8/RCShTirh4TxjrRJ7SdrulbfisNNWVLUtrItNkqLE3WPIdofFgOPT90
gNDz9aWJsn3HQ711EXkWl49aR9mSfWvDMGNenBpcCqkDXxw2mMughXxDWGpa9bSn
QWpZujMN3Gi/vBeDadWNNFfqswmg+CpOkD8jdhyzFgkE/bir6pXuyCHj0KrtrZkU
reZOoHIEaZPLct3WKnVAQfaXY/FfnUDnz4Zb36rtmTPuWUlipZv5aanMsWocZN1c
dHQEDEVmVNRrkKQurjZilZHrIPwMWpMq8OpHwtHdpS0HGCWiShuQ5GamNRM9fTw8
4z3DGXCjzWmIylh74Fpxh7QR3BICYEmFv9WtJtZARvNyuBMBzR7W3LJ2pe+eTiNW
JlikJQ0R9Gfko824jAtWIc+60ceoqj2gdzd3bYblh3G4QrBEfASVjPbZqS+maUnm
cHenwumMf8ycpei74dfyFpVGKu328GxWGePqLdjibmeNNoKcX6uHbGNF61alUapH
Sd2FOgCcsoHzdLVLs+8Aw0UpzytzGStlXzX9eNIo59/2W0s9+YG7ue/htaTJGZm8
wTFHO3CJIDJLML2g8PWbd9Fdc6LnSWs1vTm8SDzyuEq343CaQkvdoXOLwpMOKRo8
27ukivTxFCldJFciFz7EvIIb6fpk+5BWHAO5zEfTWeWnt82fDR/39rSwXuu7l4iH
TqD40Yr34igoXJWMqFsguQMkg8SU8XQJ5s2sAEW1oe4hCBTFQmk6kWT5yY+SurxQ
un0EhR8LijbltcmwT4qdzp2Q/GK99sBTaCml2LIzDr807JDund1d6iE3foNMwD6c
34+YLKOovqn385eE+Fsj7gJObXGvHqLGAesrcP+WqdoVTebcdhAAKCKB9soYc8x9
AOqFtjPTrPbTedIndZ8pbgteXFy3mVkerPDryM/tVvPxwF/aqlvvlecjxSix4j4u
cCj+gsnScox7wjvAsi0BqgeFdJxJKmFKmPEwvkDJknfFc3r+7Jl55NHJoNG6UEQL
NnZXlXe2l9Z0aq+1p5/zk5Rj3v1ikWDMbGN8HV6X98GCGBGtjBVHWlGhqbblssn3
9Qp5TWvf+JWsN2F2NAIZxVlwhqZGo/BuRvwAc81O8etKvVx5azxlTUASzE9VX6DD
SqTCgx1a3EX6qyhGy/B3xGODfR/xEe2qJnsDWjhbU4iBmv3L9OE+DJGT3AvEnT/B
owwE17m3MDUMhExBg/mMMoALXm2Q1nLu7wpd7WunA+RcYnsSbUs7o5E9vWdJqJZh
zCmwbzL6h8+t7q9d/5v+HB4PVmKmq5IycaDJ7iRSML+TIGRNE/sk6Yhs9xpGPoWy
xcbsvhpOWMtYmoj1jSlWQymYtHtS4MkLiit0FlwpH+kEvMepFf6GvjGb81PAQmfW
mPRC39Sei33DQ5kJAhr7Z3H5i0yEXpv9Iwz7Wq86L/YYoPyDd1DumsMTv/bhRrZN
oNKy1nH0hamaJZ8GNKynZH+/POJSBcLTTgcKWcNYprTd7ucG5fUNqAhDLrMnG4oa
PPJiLAOSalW6/l+ptGLdUBesWr6vHNhY7ss7DTtW1XNrW/KAihrTp3+hdtz7cNub
AiIyz7ePuXvJfGG7HaTTk+kD9sLsK05aVo6htYXiIAwN2FsFzd+eMGMSVaehniAG
Wi+oH+ai1fB1W3teJ/8bfYyJJUms9Ahuy9U/SMrjr9fBIq+pdrF6Xun4Z8fACisr
8QUa3TtKMQ6gXgliaSjyVz0xg3xYKfMBkmfhIIeRe6GW+KZLa2NslHDhnUg1BDRf
av9LO4TIsUSHXKaow3Ay7MwdNbd9tMcum+p8EGmYNyQBLrobT+/K0FscHDZ2txXI
4Q3fTYM5SXR9zyY5/kF9teywbrsunV9TbxhZ/fHbgf9IiIrlMd5NagYXg+anUZ9h
oy94kBXPN0XTMnYyC23NhphmneszTuYy5g4DUBfNrsfDyuFFis9UxT+tqIkq4Fp1
wp45ipc9UkF5IQpQyApT7MRlTtj9ZbkCv9hnlsMGEWbQy6Odu1M32sjgm0x+of2V
Bsnluc5kXPxxaas+LmYtvCxxS9LYedVPTrGZNC1fURoE1AEdEcz7VZNkA1jvu5b+
WkXCtS9ZVEfpnGR6L7lg1eFZMtSVRF7A35rFYHHHHhRVl7MBLx7/ji/GUMbu/BYR
siDhGTO4ZVYDcDw26dF/AbtCnCM+bVu/18k1y6bTu5V3mWfm+4RafhMmoKwGtxMf
xSva1hSvhHGmj6fUkpYyUR6R6HoKnQgw35TVei41b2ShQuQEs9tBIwLmCsfopDOg
pBVYLGevdjM+4fLA4XCw6lkbaHPiVLere/bNcm4rSXNPohbAOea/S+RUg+aEPdhg
SzoNwzO0JzLlFB/fp31nkrsLJJUug6ecbAHYX0K2Rft6QBgn02Lq+aFzHiSeXmGY
55je5yrFqwEG7uyhamb/shtZUdfFlie8R2ItXeMs/d/cKzGv5G0tz46sj2M7yiIT
Wys0/2rU/K5vIjafuQeZFP3t3YWPRM39vGPlyYjYYHQOODUSH0zBr8N85pplSrcG
1RTng1DCdxQoqwC7BK5+kva/Hwqttwo9ncA+mDIar+nzzjFdCCSqG/ohQviJ8HLM
mLKi39Uzkjy+4ar8ObiZ12uufn4F0pDYE5QVilroqmeJuQ8DzNm8B5tSHHDYPb8e
OQxRvuPeJljtVU0qaJLGmm6ovyuHcGjX5N0eOrMvpKsRazRl62qqyxMHkDd430Zw
TgwFKx7shGoNBGhDCFf/y5pLSkTpfWoZx1eJbMR7KV3xKPZrnrcKpxvzscW5ViYe
/a5YEPKYAtBK1rfo1LTchK7JkctEyjsgaQV4zp9IH1oYG8l1TyVZ/orK+V29/peq
wXmeYFbZAMtRCDGURwK5UtUFN4fOBQKulwZUfEoD+jLs+XlYbFHDxXB/jVicM7kg
sXqRmCgOVhL+zqgVMTs2BnUA0y8c/V6fNwhiWUny+i0fpQiTHDzQOsHoCP2fKDAx
E9rHlYznOti8pbDayqe8l3WZQcx1SyHaHhVEa1wm+o6f08UGyeVuoNHBPKlRs3MD
/yxxrXSGzO41l4+EsI3Gqi69VwG2TZfKkEa/jfRPOFGNNAtQnQFwW4A/CnVe9N5n
gthpkMsDngEu1G6CXQPpBSwAdqILQ7HQRXkTM4j+LYopMe+peBmwZXLZqMlqQmZo
Szld0ThkcJFbjP63ECFzLi1+y00cRLN0qR0jRcX39Hwxatz51SoR+7hc1WxJw/Jm
sGzBCAzNX66ESYoqSC7Mq7we3t0FhyepccZYoDyaGHQAxa1QFQZoiS5Lj/E2aeUA
Hs8Ov1WTVv4GPw8MrTPHlwuV0iqL+cgq6DJILfKEL8SGz4sklT1r5o07TegT23/4
iwgmBuNgBaQMsspqVpAVClZLJyedVxZVZxb78inpGUit3MElMQQA0dL6JrPfftx/
LzH6myaFNeRMbrvlSQLvQrHJUt4AwAPhh4hebcedOGo4SLbi81PIfl8UwsuHdmey
lNKLgA/f7waSoSP2k1BZY1rWm1xF2i+mMhWyU8ntdgywmBnD2lozoeLkavOiQ9Zq
wyatgIm+GTgi6C7b71jmzSAXLryXFOsg4cMZb4CGBq9NBtOrYHEdp68KvwzWyXt0
UKw0VZo+D8HxigdFU4FveKrpbZ5jU2qG0ldXdhhu5Dw6xhOchCPUmh9dSYC/MzKJ
G5wLVr9wCiCYIU5IXtQFd1OSl35/lvtgya+hc7gVsWBl5jFtDmXvBsGjBlVZkMTV
yPc43YeeKnK3eZy4cNj/zO2r8k3y8wra/gfDa9CeERVTEIUW1D0PwAbrgAYcdcF7
txHG0q2fHrFc0IZqKpAe8QO0SQStOdFUslRZXeYDqXXPxrc1eVw1jCjyAL76srC7
neaIidbai98uHa59w8YPnwlEoxd2iGsM+9ngirMD4p5VrQ5CQUR5UhsKcpNbW+88
UIEKO8yz53eSaGNhSz+Q91mInEnNM/8YRlWI6fLuN7lwBf0zhVXAT8g7taRgbS11
+E9+G0np2KcEQT0qh87swEGzVhmVrpsnqymNe4IfO9zJb7mSUGUP7dpTu+sQGXAh
6GYYdRuDEg01SM4iW3eEx2PDI36vs7cLQj5sQKgyLVh++oG/S7VGdbEIdLDcpQBl
KDLITnMJaoyCRKwd0bIpbo0Mr9chr/5m8eRKjvS+etopalZWhq1vhT0EcWEnAhIw
aXGY+1aEhQ3EUum5qRn7lsaGntxcVrpVdA0Pa9Vl+XAQevDeMIlvBH4Ps2nFSX5E
xL5yVZI7oa2MiqYuDBBUIQH1KWG9aqticxwoJI+R7IeEJ4tQ0COwhzxzQA20LpuS
dKAV1//hnMrB+Ja7o7PuT/8QeM4uaZ/5QdD5gmuUc6LSUXoww+0+RFUTdFrUR/s5
87zubbHbg6SItNO6VsUDyooD6PbU9Z0fCvx1DXXgr8yRuWSlFiFLN5LAaQT4Q21o
Zb2DIdvi4q3xH3bmi2LL9kGrNxA8GllB+S7a7/Oq6PYgRdCIRmANeONLfYM0gXSC
Xoqn039+arIdObKl6hF19gNGsWSRHXGuSVWcbLQ1/pyL4Cep32aCG83Q9ZRKtlVM
BKng4xJCsU/Ujtem/7f2gWTdAcmuJ2sKobuRwl/oOuLWgyxuFdcrZYGTnKPMcHnb
P+fcQtw2o/qWD3JbnQjK8l7HZg9T86UFpfxAaD2tgA8MzmzctKJtspFDvD7Tp7eE
PYSL/YHzewYr0uEPW17njkX/BUHbNgLlx0onQ2wdb4y7yB7T0SHI1Nn5bhGvb8fL
oRTKvO23aZfuX5qfqhya9hNa028P8dMMACeBWLeLTc/R0Lr1R4i4UAE16hz09jFE
T4z5kz96SOpXJZj39uAGIEKIP6tmjCqNVomA3ItpcDf66FBHP2vn8CPktTriFho0
arQZPqKIsyrP2EPFQc1eQA3tC7xSVXrqzShplHB6RLsvM9WRC8XVgtf9ueu5FciB
APvKyMKfURjRt5hk7yY4v2IZ0AZyBK+XaYVYTCBwmFTGkvQE1Ae5v5nkPIVmQKqv
+JsbT10e1iXkYPdMkU/aslJAOAiPOVkQnEZKGtAoQyKsPeAfZektbkPdbVbnLOSu
CZ+gQ+xEK1Yj6G/VAZnkncbUrZhcKycpwuIa1EPEeBHnFrslTuOhs467rX2/Glh4
d3B5FXYp62C9+avEZCkPS5VlQ3cvLGX+M2D3zz5iHYgp4Z80Kt16vo+xIJAe3oOt
bfMo1iSJRUaoOH8H96E/6SM+qSRx2wdW4QujmwECrgZ2eFLjwLeO/lAnn5U0ktXl
xSKIj+4UnGQStUPORXGk1t24UDtY3ODgraeG9v2nuHQtymjveY/K/otfSyDh/HFp
d4rCZg2WVqkBS2AyrtwW7AD+tyOxkUwXAiUmPVxTnHjj/4d3iJRWHgzZT8eJbHQC
z6q8RBSuFke3g5As9WRP70L4cS5NIJ/28lcVbmnMSUor967wQ4OxibOmTnStVYH4
1XAoZWR9H1NSTrG6buBkTG0t4XOwNp5F9wzMOKwmMQbYm3ZNNf5CZI3X4sjByXIc
PvRdb4MmK4FacpFaz5BEhxmPL+XjWdClzeforHhjaJ51TH++5u40CZqjiyZK6Gmu
oHsVsdGDNsz60fHq2CAPDrKVaP5zidkCrD6IvoWEn8PNfqaHXeAWI2OFiwcGsQ6N
5WmXXgeWwYn/+pqRwDvTRYByMSZLvZmaMdzBejdYJFxpxYwFj+RzMat9r/e7fDce
3q5RFUkxSGBlLgh7PGnMJku1gmjgdLghpowsMQrcOd+Ffp0rWRUTvD1SqdWpgG/I
ePF1MSFYhQyUSAaGPG9+dmEBHocvhqOjLJ1W2MToJ/AjQNTaJP+Y0tjgws74mVIS
T6UdEztDVbxecH42nA4HtwyPc4iMIh7jqKTNEOcWZP4uwx+hH1DamvqFINaIFDkg
RvlKSium/qVRuqrPCd9dg5LN22hZOkvApI3SYbHivqIBP4WVtJluK2GNPWcymofv
e8vLJoM5JObsW+0eVp89YLTJIzzV73tMII33GX1iX6olbXIEZVvQ2V6wdY7ZlSh9
d/eL/TpkaKc5umGDdBV3sCisklVUAPtx0mCWhuE2UnZ0bzDgLNFpbVvJny6KDLmE
NmIYE8yP9yri+Gs7JoxebD0wYtSO9h+fYyty0nRWh4AYdfYpagWDp+7WoIohyqRt
KPFK10cwKt5GWHrBX+MHjrbI4ykPIpQyQDKkbWSnpALKE8EU4sXqqvOwjKmGd02Z
iGx1mzYVWQwaZkSMrPa1GOy+kPvG9yObYonpMCl/SKbnwusXhcs85Wswog90X1dt
1ozHOOzrqxQakXclPzRugyvjY/mLty+Gtp7ho+5co8JdZVrCaHFrFHgoH/KewTE+
rySYNXWBXvHh8106TKKxMtiGdUu8Wt4Pe3dl8cVPB+2CkwZWq3srVtLSYefMOhlC
Zx1irWBzv/8oV5LEoVWAbQFOyqYCvXUNa7ecsV9EptxB5RU8wyDDuH+yc5NsRFbj
sAIpyytgcJ3p0Q/TWanwzM2g6/iYv4ZyeATyA4X70zhFFCPb6lmAeksf7ODdQAgs
tRfXsEx+Kt6GYSHLSHj8jlPwIZvV/eW5tiuEbT7FoaqrUAGkCWi5KYe4eT6MhPY3
AlRx7NqGvKvdJ4ZbIjvcRROT3F2Q6IaQjIsT2VffoalyfOOJtf4ynY5hh/vbn4aE
Xvffy4sbNPKUzMrEY91ilCOEwg6Mjwq51hjN1cWgip1oVsbNX/QTdPcKRb0Z+OSM
9tfV1yO+Lbyl3qa6Rmb9E3y3Vq7cE9CiGPf006EVGw/G+0RGcJGOcXWrc/PEIP5K
eBk4Qt7yGwYikL1sGMeDXLdUtBiE7Yg33AP5XbgKF8i6zj/h3lF0NWQNpspbDf8n
i40loGvPRwTrdjBm4Ct6RDPo/+9p5/LUO6+nRhgnX8j1XqpBTTWwpBTbZ1faeoaZ
01DtQwfKVGnUdls3IlMuOFpWUzYSOGTH9PUuG0UO4AMIKnmn6bT9KwRgQkyk28If
CrSJj4wKFKqDmpit6DKXMPOnH65OcxBEr8uhoLFcVGqSm/g23efYE2mVQh4JQFmE
Wu1gy9IxGwT07fyXUMc/aTIz376+HIZBg1UFTVqHglZcBLtK5d8MRZmcUOm+vBHX
IxevMhATyT1OHz5Rleg51LmYkZqbXVYMvlYhBjKjmz59Pgho1hZmjpU8uV+BaZfV
ZqLR3g+9QhJ2tnCoczvSLm0cURb7roKtmsTyV7m5OiWuNaQ33IVen847CIFh5b69
2ry5598x8QAwTgegiC8B72eQ8AXq5jrr5CvjgRhCCI4uDhsIv2M2OBvDL3QiL3Tg
G1pjpPhk9zMXZzjiWAb+GS47pLpa2tNdI1NcInVG7lfaU7V1ap9aMi4xt4/Yntbl
H+eHbmtmX8IjSNO8prO2or5fwYhsn+AHQyDJpqsLfPiXEX6LWj37a55qmgh7SnX9
kLVnBKPUc6BsD7QTfznsyQENDvqjL1GvnHtlhHlt/kdCLNMJE4mpdaYiOPvAvC8J
ii7h/zQRQfXuhhJHRZqeKefb3T40IwsH7KnQqr2qEKQbolMY4sU61qS89K3tVAsD
rX/coA4SgaRivw8qmyp+e8SQKR3h46LN8niPMVh8+Qof9ipMROcdBo3PwwfyemdW
2Q/NeiYsF/R7H4vvZoRKGg==
`pragma protect end_protected
