// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:35 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
K2MlLoQ+g0hA7ZxpdfkKlUUX3nWp8jArA2S1GXCfgxA7Z6H+7/pNqJLtv5MuhlI7
jUoxmyuuGWAwn7G5BefWhgqUWAgdo6MP+OvIB4rP+hyw14BSra1Qj+VJPvXi1S2m
AHyZr1UlGmmsv7SBHqHkSa3V7P0szhlhaGBGCXXBNFQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 176784)
lJJWUIhtdN/E2VHYNXxtW1atUDJ4iuRZpfD8p7/fpVnmA5CZ6qR8C4bPa1y+qo31
x+D6B4H2/EAU5XZ5OgoEroRFX/PGvrxIq/4i/Do2bz0Etz+SmpBNiS5b4cGOvz/F
m0zwEo7jx5NVPUV019Cvqy9U4x0XJTaOfeXr5VacxAqXIOPASz5pJW2UK7fgcSFp
TOUtXZ2zyKq8ACchiDohuVNfWLpng4cW7ItRtFxANLs2T6Uql2SmOQk2dWR9+paT
8LSqF+uNFspMYO7mKmChhzuE+09TFymrJUlv5akWuUQh+ZEQKhpsp02g5JqLjuOd
W8hOIjst2rrhFYnepqh3G3ZlHRPIDudyAGl+yOOj006p1ggByLY+a+bjJhbWRB1R
Nmg/ZqaIGI00krv4sfMzRgpm9VEggySFlo1Gk+Rff0r7u+XViFMpcwB9mKG31ror
Fj/XUxD5ZpHVWJ9FRVyzjK0wmaYa7nAidZiw80oupJ2XK8/71bAs1xPRSoBG5x/N
VtkqOxb0I8PKTz7FGpi14jCE8kE5Jkb6MNe59eMiElC1Nohf0fIltzs0Ir3OjOtt
Mxu38ma6PfRmNJLSxK+2ZJIZAub0tzAmxg7drTrrMcFuKOVLsZ96u2BCp6RwoC8W
YyIAxxgcfmg9oSdYXDnvlXLvUfj06AYR+BYOSQGguIAdFeNkClY4CE2qdwyFuVkL
t8J9ZuF5YX74AA3ldxjswgMdAIXMO1b1sV6sh41PrMnARQjF6K0vbLE14Fxkb74f
i4vkB4qdVqjMa9/yh4TKYFZjJFDWDZJSLCLKRcuNE+WF0H+p3KrWugNwj2HgGyX7
D5AJ1IXfd3h4L/srOSDVhPN5W9vt6CkN6QuYhbOB482ShATKBZe8nBZEoWYOysaq
n0yG+ctvLJ2kSVB1/yKGv4q4LYsxSrZGqJsql/uAotclEel4HqnHd1hP8tlgg02U
E4qYGVJ42fY8E8XzxwvyitXCpHnXSE1OtLc2OfhyGB5INNktiBfwiJbCVpg0aw/p
nCoEhQLL/CFTzsCL/E8UJxYVEikCMQ1aXc+Hsmtn6+/KUTDauZacX22wpJW7bWnD
+bRbT7U+CUzFBShMCVCuh/iFc7TpOPBo+4bLmUrN0hBIWPLMnQvTArvXsAgTbPz5
jqN86Cx6ljW0/D1MAQPNchfHzY1OcRjpKloMcZ6wPC3p88stN8w6pq3aHYTK0XL5
d2rMgUb34pCaDGLKafgJrue8k/rcLdLsenUcmpFg+KX9KXqJqo9Gvl7Yrfbkv20/
81EAq9+cKRCF9oR+n/JPeU4/gbR44nmQdQeDfGLjoIr0S5ffIK6GHPMWouBuSpo1
rfTlR43n8JWkJEg24Y9AjmLhhXJp+J5Sbeac9J0FMPGthjrk2Lvz5kfdz3WbY33y
gmU4e+1Hsi7P+/Uu0UMrrLVKJ9BMn06yje9uFdT84XTxKRFCrgq4qhSGwtIdA6Nf
SbASMW/ZxML/J5aIvh0lgVgH+knl3HzJmMG/ogeV7D6xDuwZ7bUU0btL11R8hD71
lpWbfUPYVVOyhEhdjLwBCXomcycJ8M9JQ1sVLmuOJRxrHvVYKskP9SD3tSdqfPS9
/vqsbqwlNhArbLFMJOKD2hce0q/rKf89UIlnmXG1cjM1RP3IxqSTOCxcL6UzbqV0
OQtPkoqqRZfdcB43i9xzQvhRfpJkFx9K37NJWFTEJ189GPStadX98E9vtFW0cLzx
i4FE8sWTDJ3fRHrpVLqaRMUk9PaVeujr6NY748KST7P7zFiwW2YoaiYEkvItmAtw
BjXGilUyS+3lWsWcAxe6Z2UgUh2x1Q9tj8+Xn2IUK63nXyoSDhvs2jLOGsJokOVS
60nUK0TSSntblr3o4UmvYFNupJv1Ok78M/1MrXPB94T9kyU9Lr6cCIHit4i2xtHp
89HPUCPKsaEvlVvlKA9Vbsq/WRDamHZbTd9GJ4xrxVVAXvEFWg4ZSEZPrOaQlJkO
Jsr7HnlfdsLbDmcA8XJLv1p5vJLtmH+9xL6phBRLVVCsiNESSriHqmOtD47qPvGp
3Jvuybx0mdQ8xGN4t5C5FWh+3nSiyin8XwUDedgjci3g6/SKaQgz8i+ea7w4X4P/
3RxJVUVjnJil4MnkSKFZl1hCaQhHo9SMzq3HZd2FEzKtGYouZqMFRgLGbtp1SVQA
YHHNjEk7oq3xyDRtJu+li+X4Ujsx0pkwkvmgWq0pvBHzZPRwqnuUMiwwDyGe6ufJ
vwe0vqdAFZ7Cy1AF+QoukxeT1yTFfkcCYWmSWGXzGmu62jfyNoIdnKYtzYmA1CmA
Yq1yJpnUjh+4MtHnRd1qtY6djStM6oG7GitrUS74Aw/DCWmPaF0os0UcJdyBePaB
58uUeBUQK6GovAKQL0FWkixXZgip0j2t3QVuL2IM+XvF2jo/9QpRWBa/UFyrnD7c
OmDgI325O16fO8GzK35JffZQ1DjtDa/0MAo6Y6kP3yyrFBBW+REQpYpFGe5fTX/5
eRc5A7gOk4/uApZSAcKLWok3Bj5W0UO12xRWsY5rXE0iRf/T8yocDkWa90gwP9BT
3OrVVNiTeBSfEBYwyiCYcZEY5/u5ZCy3pu7V4yH79nadDlpl6Baco5Tyv+q1Yrj3
ZGJn8cbfcS96R0y53DMobmdz8IJPl52X0V7NAHw2BANygPEtqHwAFhJ6tPP/d+RA
/X4OOfLH3soHLbuqZQHaQE1Mx2Zyzc7pW17lFSBo9/JV9OOtuJXqEWB5E4/92M0Y
GN5eDhsbADTwCGuKZrQJ61l+eyysSz/LOsKCcH0jJFw4q2io607OM9+0JvmUyrLm
V2SNt2QPxeQaM3ITnLnBgFr1/J2hT/Rpwj0EmH7izHjWN7dc5noLdRl7ii0mIWsz
ixjfLRq0EL+9aoS55dYuwlgqmMcXK3kSXinsSQOVZDM8aVT8COA8Qgm6E+sBHo2K
F5+RnOzWWpVkvA0KEmdmacnawKMpTbfk0kcPIXSiO6aS74BBk4orX4UcCtwnqVWg
eOeqbgSx/OefBC6G/CvWWMtA/zBRXZka9o8hdg7D3r01MeRSgl6CL96BOqeAHUmZ
gU6+zcCGSsQQMV5Ed+ZYRUnfuwsF1nTpa2jnFc6J8kNJaIj9jWjgahbagHi3Frfz
IMHLCfTjIajHToaV0O7POS+uceJz3mRyB37mRq6wTezBhnvPe/SRYbPzcpxBhNyN
QP6nHVUno4T0PAUPP5683igfOGIDgpdBy8ottjfBgDsM8gcKD6SH0tFDnXY3MhaU
mfprg2C4Vl/W2zqja7iwWrfew/D4nj6S3YLB0IWwbYrO7m3xItt/TUNMYRjhQgpa
mHmLVVPvEjFA0hRBVdngI4hhgU2bFiVkvLmDV18ZjynG7OgcX8oU3kyB4jZ5Ulxm
8oJN0d03Jf3AIZM4A8w6LrVMtNnvSzwIiGw0AoyatYqvo+cExwXdjEdadbu6PZdg
X3UoFaZfstNovc5wlYGobjSygIDI0Y4+UBvmS7aLt4uDYMhWE113xGbg0NWnD/12
AzeM9a7JGXUR9GdQO0NErWf/0Qk6U/qKwk2PW+HyRz0OGl9OrGIOAWBbimAW8VnJ
iVcz480MCoh57kzUh3C3i/+YMaXPQ/lFvk9d55B19qk63fsd6sc4nM5fQkg5WNDn
zq3mv2ptC/tflsg8q8RIN4O7qO+cko084j05Hkr4nlWKxuY0rBXCxge+NJIV+rpt
YYMX8ctMjMBmGs2QnJ6Y+/Wn8J3HCU3ErDqoLNo1Ol5bqFyJelqAgHO6swTH0I7M
0lKw36+9fYFdNKG43e5cxEuHWSl7zFP/aGS6MElWmIdncwHMiZDd7SZn4jKF0tib
Gj7PqYItH+IQefDFztkzIXE2ak2FbwG1LwBy/E95oD+8PQV+7a9BDLuLN0GBWMH4
XAFv+405zOC01dAfk+Wvk7A4RzTaAKx4dJ4Lcfco8w2vRQCl1+xACEPpi67VxhGO
v5RyXFSzjmk61TlpIoF0/x+awLTeae3jjIvJ8DOrqWM9RsccmMSIvZOBLeooiSh1
N9lFDVEt/6i3PGvzjq0HSbHWK1JS5mBRqaJlm+UmRPOHwuKWDUun7dauOTF5H7u7
yhNRDTalasjkhLjYox0S4FbRjw7Au/SDxKojtQYFd4nzPP5OMqkRsSjIWTkjVi9O
iV5EqsG7q3U10rb8r2H1+AXzS/ThitLMjU2/8nfG43ZNRxfO2U8He5qlLlI3gMJU
KvT3Jsz9xrrOlNWgfgAL14I171gMAaJVAG48wuQjzwGeQH4QVparCtmlEoKYRVeW
X0NqvwHtHs7oGmpOWThgikvZn8CCdpIDRoOQJDj5zJE+BUhuTCcVv9l21iQO3GzH
LtLTkrD84/mAtyZ/XyckTkOyU+lhxV076OSliDBWaAP8x48tOF1IOUJrSWzXniaZ
/86jhdggQ7friqN5RRwKWG0cs+IGTBsOQzdJQH7KVKCvvfTjoBdsivkWRX86lITj
lGuKqtgWTu54fMscoNysokxXSZTIxAq4DLc4Z+t9K62uwQFnDaOjR4kFuheZojF1
kUW/Q0P0N3Cti5dLUDe6JzVRS7yVs4ZWx34xv6yJkIsooUr9eTRg+ATAISNkcBHM
iyAeO/mE6GOooluDcHn2uLpfbO+yMHYLhBCPjxrGWOOzydJ+dZv4YfnUBr4Gq7Dh
2yZczHH7HAWo+eHrkpO565seislmipM+RFmYWsHD2+i+rdjk1Tcx2QV0FdB9QfOK
E/AdA0X7Vi5P0/d453iU2WYvIopW/+kczvCbO+0RPzsI0imvfusveT+2MGbOJWmZ
XoVnXM97x4sqKabStdVLc4ltz87zYD9ujixJW4ONZFWSeeTJWJg72xAqdFG4krR4
8Z8knJ0HIaRm68Kv7wklWa3eRN+buhuqt5VrEMS9SxTtqsDzEw7Pu6PRe91G0rf0
GUMrbZhrOz1czgfWD/sMQrlnXpff/i5gFmpc3wPP1MnUnV6VnF4AfgX18illa4XQ
zyJDFJDA21r6wqjhKzKYkSIY/fxFzBti+zeU5mdbwocMX7vnMeIUXKkL3r3/xUVt
EtqF1SD3nvn0uzZUpWDSpJ4mX3ISf4o9EH8gpkVtlyBE2cn8Gi25aSeWa/EHLGgY
/3SsycK0hebY1OTyoPKmpf3xXVmjRTHlTVtb2NpTnxgufoZXg+engdMuXyhGlfx5
jN740Ixgi10svAno+qkvtNKT25g0ITSZfmQkP98waNH3kQBN/GlzCSocqusWzPAX
q9fdx5gCTzsqDiyqWKr1qdCX+uHEgNC8EIsq7vd5fyFExpAWA3piXq9h+t6qJ0e+
cmTrPlQgdNLB744LIwqT4hEImdMOiw2KmY2blP8uPmAtw4MbaNn1rvFMA6vYPNA3
Yyo12QuS+0MgmjQrxGml6XtEOi90rqRA65yKfqhzSfCUE7LZ3iyVyiUZNnQtSuvX
GobtNhOeiLkn2GLfjDvxYs2tgfhJ6r/IHiVeJsQVGZ412Wged7hLjWzp1tu9+gkG
9OGgvSNH6UOT1Pb6biGdBJxoUapZ2ggM9x6KgEmXlhrpFXV0Lcq4V8/2XDmRzTqe
NZFq8uQMYB/uWdo1joyAZ5CJqYfRbDq4yd57C5UrFn5dh2QTkwhUOA87lqde9n+U
RNLyKK7e/44jH85dXMtS+TEDoMvQJVURtStIrRn/EyqnPRbTPpsM5E1MjsyNG0TA
FP1PjXN/yLaPQMpkV39akMgFNDMAE9a9si8EBZDQkpoF1q//E7SGD3kkEQodLKm7
s5yB114kqHzl6H0yShj0KyF1bMR8RN2Xhj0WOLRHhbEiIrlMSBy7lIFo6rXcFg6n
1w/LIz08D/vfMC9aKwyiX8h+sVl0/qr5tX9MWwMPX2HbPAT7J4RQr5wXifUf+46R
nhYZMC8uwhNMsRCn2mhG9qZ07EVQMhHEIOx0ogrA9Icfz1NDfotUU8qIFRcdZ1eD
bgGXjiFanS8PhQvWpiHmu2n6m0Ywq+mv+vyBXo6M5QHPXQ/FaPQeHx//jjnqzUjl
GwBzZY748UBQbmhWd4PMnCg+/vGP0Yp4WSIfi31ypqIf4PC4dMdBCPJX5MEcFoqv
+vJh6UHZKuyzQJbZgPri75wj3noaumtpnpfTWXFMx2AEP4iiULD5b/Jk+6bANTG3
UAGRlb9wZX9SnsYiHnvHHrqofunwrQzIOrML0XzN80OsO0axWJyY7nv97Svm2xnr
s2e5tY0KsMbGJcO8jrTMfkQA1CoTl+E53be8TFZpTsA2JgumGywBHDdRiYe70zzR
kM8NIoLkNS3BQRY2cNxQg+cukRzPqhGLdnkV+IvcI0CD4kyxFTbVKy4/k+zyDRuk
vJrwpvCBmxGwQPtbuVp3EV8UDYSduGGNofN6sWNdP2oBk1e/btoxXH161Z/WABjC
shNncJy+3VjuaXzkM2g2Dwdx4XtMDVHdLEkjTElOElfhgQxWztBpLsHE6W9z4NhM
UHMrVDjopEwsED3C2VEl+iUmf3HC600oUOW98pUibhBQBUNYX2Dtb/fpusLtPSG/
DP37zxTjQhNlPFrl56vWW6/DKpqmo+AztnIE788JQnxef75MhpAiyWLBBwGTwthi
3JoqLhYyCjdL70zQAJbouc0zUaVrWiiZQjLK9jEohVr0TDlSH8OapSewt2TEl8sv
XdjKn2gpcF2t9DqPHJsFUoseQ2XPiP4B92OmgnCJ/a/7n5nJojOpk4slTGovsVGl
dN6RwtgHMDZI4nSHrxQwnt1HPIX/U0fUBa+mT0owODjjp1veQQivwrbMwIFpzOEY
vsQVYU6e0gKA7uSkdaiox4HytMaHmTKyO7ysaAmF03wPie3wGk4VnAbHN1I/UHfq
wPB2kzrLvaQ8y8hzsC1uxGctcBMoLUwUH77Tw6OnWXXzGxPP/u1lPGK3EF2joo+D
gwZhIFff825z6RaybvDkcHN5LaEuVBe8AAjFKF9rx0utxAgA+KFTWD2Ad+PodAPI
z5wzCoDglCU9VuTE9O4RiOKnZDe6aTSnwImyeOCvLMhNq1DAUkz1MMhaUZVvHple
563QJFZTe/oSOAa4ezN7S6Y3PY37w8XIbe6bhVe7zdx4sXekckhks8W6nRP1k2jE
1rx2jJJOqmqpxuMzfx3Xph+FLFca66tV9Eaqe5lmqA4+xj30GVYBgNrQHp4Xg+dW
n6LxW8ATQOBtwZ/pPESo/wf0hYnzKPxMnRD+qHpqMcAbkpDK1tzSsu7D/kBOCOlh
rHZrBBFeUqSIdqoNQGRyqGhEf9P2MCLADd5gZmAWbTMBMH7pNf3jPxPY/xariFFf
QfgYBqo/l+/J9Y8ZfQJm866q61R7R6+/ZFY+PFpeXfTGyxcOfXVWKYg0Dh3zEFtR
tUxK9OM+nqAUuT75yJP1C0k9CfgIc/4ZOrQoMH106c5OAVBxVNxQM2VbCbneGboa
RmwlQaOmlOYhP4PcGFVjZNDqOlaAKi18JTjZEYnMGfYydHQMVh4b/guEqm85+Ry0
BOHk03VhYUQfyZ0jMFlsU2qHCpJvbkj1W3P/6su5UAT9so3N/a6CQWL19RXcLcd2
K1asCOkO8MtgVpjAcwm4dfUG39+ojpU6pwGvsp/7oppSlpGzS5rbGxVE7p4GS4gH
kxroaPzoQ9HSHVwYNtLxdQrJoIPPkjbxG5ldBo4E1d29VMWOgtrkp3LkmBD2e0yj
6BGP27dUnyqT9wIndqfGhYDhdXYnRtQ8JGaVtAK/5tp018P4Goud8rGkiMrap+yC
Ijy/hhbE0JOc/3/HyjrmFE5pW26/+SOc345NREbBqoXGBeKc48khO6fZ8+FSC4ko
SVQlmRg2dUaYhhR2Hnx4P9+o6swmb06IulY2XvNGvs6YPYarbDzm+x3Oyw6vAPX1
W5+CBXgPbI+axIXkOwmraqMY+ihYArXfV+g1xLfDdEokn/sEEhSNhlo68socWl9V
mJv/gb5UfVWD0F9MrTGDrKpYtNRAhHN9hU683FUR0jNYb2azUMCTSYZt27PQZYvs
vBvsWa0d5gujPQCIJ73r8rRkALcn160ji3TEMvLXe9y8lanmTGH2j1J6xVkpvxVf
YIPGF8b7liXzhwBk2Ss9TRYO8KiIR0UphgNzT+XgMR4BsXmCqmKGQURZ+/eZA0+m
BFvZXVLo86oFI5cIMgjmmJR3eQGKPPYJ8utVOWPc3cChbXqexqnAhzPBv4muS0p9
VsQC8RmR2ZQVcONAHdW16kxdNe6xV4komecd+R1YOYOoF6XwtPdtU9Wsf/BLSFDq
n4IFfo7+u1nQhcROG6WgfM01qqJyuRok/qsOknaHw6hSqJOYslT3hw+NU8xYwjKH
fPg9R4VuYwD13i4oZLcHhIgueyf6EFbEhtLXYuF9D6qRIqT2IXQCiJL1dG/j58VU
DIl3OQ5zIYB8yxMwDMEMEE9l1m+FBjMt1LYY0JKqapEZiYKg2y09/UwmMM13Cegd
7WqC1WDzgwafoMHZYMFhkMs08ETUexI4K1JbUSnWOAlOBg9/G/+Wfw1F4k5GHcXf
SNnciI26dOAGYw36x6knO4ufZhHX2FSVvT7LgESt7Drcqm0Z3uZVLWmNIehbta6q
4xCaJvkinCMSXK4UiYS1obkISIYj5Dmafd80RzD07mY3wvpMhrXGpWyuG5zpOhpS
uFrc9lJfOmQFJgGBl4h2LzhqP0eHLSsS1QM29MCgHbF9wnF9zcy+Jnw8OjSC8HTy
cqH7EpjZKycGmBRwUFhz17l1mA6fCX4BM6ipOYrWvPjOFwxyk+CgWAdDROhq83la
g64lytPtOGQQKIOh208DiyRSXxZE6KYP1GsBNI0NySuLfHkfQpTXDC2LR3/85My/
34BzDCrSb09WOU0ImnEto3b1Wb2F51nLDQsui4sp01AgpvSAgFI0CjM2UgLNYc9Z
XOjatM4h4Jl17gI93ji7O2e2fb0lnBPdmML796DdPHFj363pGaFW53v5SKNGFI6I
I4Lzmwe1Zgxo9D1RC3Vt5mCFclarZBQpcHv7hbFRQLThlMH2pn1iv02irdITR0Dc
7/q5uX6ANgbbaJk0PR8ZTa1Bg4E89gxszB0N3NHctR2DDGRcn/PUe81KcmYvenor
4znMKrfYSI3rDwrPI2jY7Tnn2Qg2nmXEvVKNiY9nUFStoqaGh7sDoUutbFrbzj02
73xq8zDjLVRuxu23wgj8s6/ePC6kvHCt/ryh/fuO8j+7xVNit3KUPgGFKcqLXUe7
4W2gJVVYmzK9hCY08LSbqcWxjScsnN3xeb7qcH72kf7onYxzQeesjn48SCeFby7j
Rg+bY5DWJGHUVwlse9W2ALp/vWYuIzjE5eyFTpnNNp1ZA3EdaqLvAOxGAgp0r/BD
GCQX+9ewmmvgTC4RPXRcJHQBWNa8P89YogyFf3lQqtAqPXnsqDqePIcUvwP9cDEJ
Txyvrg5penQQb58vItDoUOy3wYQkNXN15y2d1oQZOjMR0dA28MG3IKn3ybFcg++7
D18dT0DCZSyVg3hf6/BDG1a7VKB7cY46H93WX1M3tisA4cNQR2QhwujHREbga4bU
ukiGs5JgQHwoFhjiHf8lSmVEFkOsBtco5inYie1D3r7cmrdC67v55IC68zgPNdid
zdhRW0+2hY6GHTKothPxjG0MvmewZcmumNaN5oRUVu2uYD+kCK5AlwTpvVD3HVT2
A/P/Nssa9z6sz5t2l/YENqMldGL1V1jZkY70idaIKCKLWC1yWtEG+hAOXp1Vh6D0
jX8AedAwDNUpvCIR5AFl3DJZE+j+n74jM7RmbjjjUxFWdtq7P+9wzDWzWk82qV2Y
8m4ai783Y467cCgoda7yDUXWHr3zXGnZF0bHEhebzn6OGhOB9yvIwMaNLmI0w3HP
5PEgQFTSW6s7HkrPpSVa8d0bcFkhSGOOfgnlRUnwyKWTmafiDoFJDXb3mtHYqHdm
y5PwgF12Cm9th4RAhBdB8olMKecITUA+rtUMaGpkjnklVmUQ4vWs1HSkWoi4eD9O
txw82XlWvFLtF3x7pPnVLGCnCVN4Pbk/Z5nZwgNm8hYykZI/EZkl5nPQp62noNnA
mZNsrNSh/7kgU361bt78zg5L2WiRjdu3PgjLSUzH8jI3YB4S5pAoEJVbgjy5QyR5
hKidnvMlQEhablllf885HdguIKTDaiKia3XQynR0CeQExyJ+FZZx0KaWKrVjlKjd
PYKeV5gBdz0Knf+l6On1g2o8LJ3hhg8zJRs+8LORWgY56w2qlgRA6pQcuU3ZzG57
Ro2UNVtZgpv008QZfjjOJikN14RI/uTUMlEPIqvNMSLXXeEK3GkLtk4dHaPk3eHc
ZZxNJAc8yEfZsPw6X4r6AJ8EE+6oEK6puWBWFhujTpO5Q2u6IYk+FuWUbJnM6dRt
NONaXbi9DzkwnfZOtVFaI1xaq7EiqMLBM0pKurgFaik8ERog9f28Nu3ZUsjqpKWA
j6D1pOv8lQs3SvEz4mOrUUWODWuWizQt/RV5TpqB3x8ICYnALLRj7V0AUtPytVtH
boT2+ZQV3HcahCjMsZrZjVb0HrppGD5VcnpWZCbTSge/yNjqYIBsiL5sHyMP43vu
3NqnPfcsnEoJtp149l4ly6UVCzyMj7laa9QnCyQSnRkWnEdHJgSrnAT+uyWm2QrB
iM7yn398kfafz7yACpYII+zpWGYhniocfXg9IWys8JBjePD7wDNogoFMK95ob0DD
9o1DwzyHTsxVGytZcWZE6Y0didgi9ocGuj085ZFAzlF7u441lNvJryiyWgEaT9gE
Y4kIQTY3vMLZHeDw0qp776aaCsVhIebMQWJwC6aD4UJ4ojt88BDCIKttIutkZb40
fz2gT+WR+F8Hzt3VEu4X+/5EThhZ6nQ8tsvvvibvr1Q7E5cWKYzhplmoMXfmuWlB
Ak7/AeCC9m6GvRRBTIaMMU5f36ICATP9dWwWHN5cG1NCQTDDHoB9VpY4z38hVhmc
SkGmV4uPZ2bUkXMQz4uYxoaNAzm2YrqRAmA1WHHcw3niKodG2lAwJ08TroirNkWb
5A+FXm4Uv+3PI8wvbWGD8ued+jBiW6w8JRZrPXto0HbgpgCv/1mY635pnYTHFonT
27pDLgDg7jD98kGcNVfvQRg6F8gHRvRbOF+gIvOx2KjYixy0OCwRptRBz3Jr8hPO
9AMBwx91398UGWcZ8DD3IQ00DTMUSAL1fr9OyLrBAw2poztmn4ae/hJmCmTfFfww
LFTtNkaX0HyybVV9n/R5VQ2y/oAf7qISUVQ9YVWbU1yoHj+B68f0b5lKc/1hf9W8
7bF1e5gOfpIRRII2AbMzSH+AfHT5A9Fv/uDeEoxKcyZxMOEwd8R7hhWM5KMQZySB
znPaJB9VQbHtV/tDdbCGnSDPe8FV7Iugdka5dlSsv1n+1xFT+RF3TWaVV6kcS0hI
EVxFWd8Ssmb8Zbf1MFus0v4d9hm76XZByMj8WHvgtAyux595fNHOYcphl46rmz+W
Ofn8CY8wy4jOfprh36g1aCSW+1wkvwNSFAczRM29SUXJL8Nw/h4rvD//2bP/lfBf
N98oJtOaZSf4efX1tIRgwwvtRK98BGlzbmmOPLGJYo5ANuLU3UOHyNngb93zzbEo
6QIZJXuZa1InpkfM8g96h7djCbDYI2l3u5wNYXqd3CG/7mcxkf8KJsGYeNwqEpRH
YFgy5/4DwbyltsFIH7teoavODqB4NDAKDIr1RGoUnqsH1Gbm3hYp2wocPJvNOBIg
aEqoqTxosy+h8Zj3vQ1kih0PwsdpHqKFfWUlSuymyWUA1crWgfhlSK1JSup0uK9O
ugHMr0hzfFmgHg7iB6d9FcrNiJ3e7nV2gmnyWCgOHKGHTP0yj6tqyuIWjon3cwKw
6RTP0vqc1uu8GC0g3ktIyQkxL8+s+/nqJO3Oel0T7xsH8E5zfTU4lXFZr21aGP0v
UV9gCSN1vjR97+8NgcuS/cFDw2QojRgu6rIdVBy2GHuGCIC/JiQQ4GNpjTU07iw1
hJRN1gVVBQHlmXkdp4Vpvu0urlNBz+WjBgLbfDrUJEiXLtqR22iiFpSGOWGkM5YQ
7uKnq3iocAPR3DPZ3ITywPp1Cj0ZwFnC9FOJUFQTaM5pAQ/+7MwYPje6IYzaa1kC
DXu/5qdCE98xh0M9tv4w0GTjj6uostcqkfijSmZ7gGfe8Pfxfcc4Zcyhwhm7Fqqe
1nqcrFs8Z+DkteWmMbXGi8i0rqqyPJ/qgqw9tq2KFNjH+3eVz8rgKFYPDuXbqWBr
oBwlN5hHwGXTsQPaPsnE3G9LWwLRIEYg3+C3/wFHu3tME6CbrEkORVUaxDvkOIsM
GcDpBNWmPuCkJ/udOGm3BGjlXfx2pmMKivcm9OVXifr3oLeMi14h9YFx4cWZG+L4
ZeR33SaHYdrEFkJoTfQiyxkeFO88KKkFyZEHOcs68OSFyHy4H3M9d9SdHrPNLpXf
9WSrrV/vkdhw57DLihISchx3UZN68Vm5LjHaD7/BA0Zb7QaXsSwHsHd437UPVR+z
GZzQhXaWvFAEuhlo39WhZ3ea5fQMWCWe1pGIg+0n3nDEjVJ3qryVkGa0aQoG+wBJ
yPYKLWDi5sRAEEG03J2xv8YKgzLlicKaTAUiUdynCZDTJRZvWRcXAInSInDyNQV+
w4zwhBNMIRHEBYzs8p8HioznQsW/HS2XE90ce4ZzLdd88Orbij9adRFvLGoQcAEQ
bmSsICg2U3rgNPpQwFa0HCI8eS7gAjRlv3yu5t/5xnxAnvWiQuCi5ygbxsqijXCz
DvDF0Af1GajWUfMNwFwdO28so7CoGSYFxvbWX1xy5AhtwdTPLkUkaLaD0Mn5ls1Y
TlxgPLMet9iDUyd+G4be5XnERZNepnHqcJizLuIuadoP8cizk2dhz5/TkCTVNXdV
mL128wVBrweCtVRx/ZvOV5x3VaL+sq0x3roZ9BjMIUfbmujliydkyf/zUvBFMQc9
s7HI/RypfxOv7OKDxxW7fsYTm2b6p8E5CQ2+G1LkDvaccXHZ0kEhUxHofh/Z8iwV
mbHTEyn+o4aDJJMEwvX5b0fUrBEb/Qbvo2sFASrgc+yi8tpOVlaVmhHElRe7lRio
oV5OKi5J5cYoEewwLqcvtFGjBsSPY8WMFicElFo+j+uogJYFK2v/d1G9PG0YsdUj
vIuhLgyX7nrvT2xSkZnFUCOxVugItHouH2VYuwa9qqyv5XvcyEAE41jIBOjEnJbj
b4hg5po9zwzwECKewedxmrXx1sd6A6W0M2zjR456dZtOGgp1ibcX91DLW4jMyu8m
x9YlWzE4qXKr9suRbCGtHARJZzl77qvn64MYPc3PBGl4/60q43LcHbKq7bBRijsB
1odiEEz8V17r18MIQAYr6fHPmmfLxmVg0h8OqpBjplH/eVVz3dc48YqPVtS2eXe5
Kg/j6kcpKGlPnbyZzaEBnV32c2eU8RmcI3Nuv2RiaJguKjQGOOgTkTFSRDanMaWQ
74zs2tRbGswunishn2L9lAtx0rGE9iG2ZliPtBPgnXsxZsWD6t1mGvk11/PApgXK
m2h7dOdw1P9rmoQskjHcRmV+cGvihTrOQGMrvgXPBDhBAuXYnFaID/5a7Hd7aIfA
0mRp2kzLWyQ0OPrOqVIkups+mQDzcRqE8C8+KGoDiuik25j1JBmL6FcISmYF+oVR
v07lmGh8YD66fZWsenhBVxASBuGLgtoVGVmVIxR9w4AhvOsvtKo9vWydksByDx7C
I1+QVygDboKe1pp1jmI443ta3MxXqEulmjxVnqFi8T1yPFM68NB1g6i3m0+Vb+m8
XVoAU8wPse9zzVki7acVG31VU7+7MfBGYeKKy/D9knzGABFbQtCxYZOMdrkRw5qQ
o/2SIbAzHLSU8imH5q5kumFN11GgCtxluk3BzGzIQ7YmEXelOPHDPKr0yizZYQ0r
dkomnntFLW8YLm+whzzkg01hMJaDVAhO7wf1qtl1zPUhIIOakC3t22w5qgTpkazQ
3cARJV7SVh7dMUE9N3Q2YdJ917kJfb6sDGNbk/RibFk5IeOgF/HVUCVBDjo0whcy
ePxY1roApyZPbRQ1NnjMTyKEYdGnbH/4h7dVQFDOyNlvpI/m8D3daJnp4Jl1ABJ1
JpocGJleeHY2OheZ0BYQ2sky7LdluuiHu2dYE21XtiatxagfNs/UJT+Mwtq7rI52
k45mgKmaBPMYmwDBUb1INw7C9ZOW4K3oHSHS+W0ckxX0DzYYbpKbpbmOBD8dxUI2
G2x4OAFhg1CIQ2zoAHOPzOrpNMfkXYJ3HKT8ZVPMU7j367ji1IeIvdJiSgGdBFuR
P7dZRuf8kgyYs8s4xVUU9lGCj1uwHwMbTfguXJK/sDdZGKzefQdvNnUrtLOiM5Kk
QlfsTqUH3/nsH2KG1B6uCrq9YVeok7hFJ9HyxKevBlBKevejZpVlFlH4Pr3Wkrkv
MicKwiQyZTLGJtnLEt9dZ2gG6/57YDRrGqt7f2hK0UIquGRLDSdVKQ5W8U2BpClq
QVJSa/eJ5brdgpLDlANR0DnqYN+5cH4wGRz0dMCMxX+KLHOtxBVen/xHMAeEa/LY
3Opmm5QtC7VkffNylCJ/1MGCNHxATo/zZIZ8tXakVbbZtd2X4f2NkQXtC8GAhUwC
qqroyLPxZJQebH70Qf+cu2rh0I5Ii7UAM8SY+239UiJJu9ceydco876CrE0Ojf7Z
5Q6tNS632/gpJgnPriNHvT3S5+zQbDbp8KfubBIIBZj9L6LGbR+PFRY0PBLerdH8
/fXMVEzJ5G518LBrcZ5ktd+Rg3PmN2jfKxRGHYzAcbtaadKvQ7cB77tYMIWSoOPb
8OLqxQo+n+RqlzL2aWPin/wp/36VsQJqhRU6flEup55OtY6j9Jgh7QXM2lBB0Y0J
uiZyboeYzAOoAaWeyhwPrylncWlFfENWGIfMkabS7eV5Kgn9VSjCvQaqPIcSjIUA
OotQCL8L2PgsSOWxkLpqDfKpAgeC8V7t2zc7aeF2GC48vlY8GqAOCDOG7PTAXLue
xg4Vj01ph8EsJYpWWs8skACZKnxSeM1b1j7Ao13yUL1MxhU6B3/Th0uI5MB77r4x
yMbYpA2JgQATqDbtrNmmjquwyMG+ie/BOWcuVf83cYwVrEvvcTznK0BcPetippLx
B7Qo5NInJjZTG6Q1gHa+Wb6ELdtp9aJgUyGYMkrU7hcSzUuzhBdVI6x0vDILHEUu
9KuoAN98cIHrF6enD/QEoyaHnC7luIL4XEYFxgUOKReN7m6HG22U8wqR5y1rlds2
62hIqlqEV2geS1bRIYIhw9icgt4ufBLR5K7DC5yIXtjg2jmveSczDme8fM7OBFL5
I7XyvkNGsln5ZKH+9LF4YcTln8bA2myJGVRpJtFDAoH+5LawPuTE7efTsJrl0oo1
6vH/l11/fWkPatzoi6UBeacPz3t0KpDcM6xScigVe4p0g6gURRpuzeYau2mIXarP
wA7v41FDLLdFRk7APWIGoQgR9JTF4SZNVP9SKaVVj88sYZ1REAuisZblytIe/PmF
qwO/CHCJt5cyFkKksWXWPvc0Pg0sBfHjGLXc50hbZiCtDbY0C0bQJ/4411aJ0I7q
dcAx8raqY6tDMGlVo+MsuHf93IM9/OC+n6bjdx6UTN6mTLcvmgbyT8b8VNmB1SiH
A5hxQioUEguvNGRbr5VwfHzcrzQFOwzAibfBWsJNX0MHeB3aJqxA53eEhhnLh0ge
5H2vc7NrmiVjFJmHH38ULZF8SCUVV8FPZvs4ZhfSnFwoj6xzYsJgI8A8RKVzjC2Z
i8vjaNT6IIgQSdf5bXYiNXYcUqUpCnWG1CMvRIkMU0o3CZnHgQQ9ekIEqqa3R/cq
bU+2etk6eiL3Ph+KL+yL8Ar4p/lhsPxakJ4v942DqdU7aTp9nrLEfg4BOCOHOeJB
HY16gmmU9ynuax1Y+yAZC/mdYHa/ROf86xMC7I3mLUAZ/B0Cof1A4rlWEkQzD5JX
xDxNZp34fg6AXWxxXvxdvV2kWg5bAONarIOceZWvTy/zEFiXExcBCZukzuBdNED1
iaIrjUEAL2nDAwMrhMGnoffHvd2lYYmKp9NQyPSoNFTCdh505xPLNjOaopu793hk
//oG5QfL7rXhoq3yrmcxpH4ghcQCw8ftruRYRf6SWlTsnNsphwH1kn/tp3HhqNKZ
rdSwbIC+AgUPcp5uuPewt99Ug81MH/CRWjI7XtivEeKqa4HgudkZ/ifMYBMG5oZi
D+8HUJEjJpvRmYhROSdLWk915BcHvd0F+O8mm5+VtdE9twU4XUw6vgCQFPHp5Ba2
Ma7xE+vSWLt8JWp3nuq4zMeFIcl66DBl4XQNRQMA7OLtDY6zIf4+FaDp3G1ZGK6s
aupHxV6ak2/dwjiI8rv3NJe/nfW8mQYSHCv6ZB6JucDOMyglYCNdhAyoGZWEeAjT
LUD+zWYtKaGL6G/ZRkUS3/JpzwmkuRPd2qoJ7QstZJGkPr9jqc9FCd2jHY0tKfnx
btiU/u7s4iAU02i/A2LYMHEHOhJ4B2FY4PaQ5hmpk09yAEiAG29JCNXiZClmLR45
z4kq0HrcjCNUsPAjvTRualB7a232RnaaOvjV6gt/H83S4JmK2pHMFQYFHSLJAuki
eCe497ARFBE0foiuXA266Yafn+cv7VhCX728qDGV5TSyjb8QTAel6gAbpVHvwbom
uox6/0pQtaHczRtE5slPVeK1VfPUoU5T3Bh7HHjDlD5dDgP/+DcI+VFlQ7/Zb+Lv
OolicpV/rfP1/cb1o9rFkQsVU7J1537vuAuBXURlOMlfh/3vCnz+DbXay3gDcuOx
17u0AYDOKG9tDxlGncTeWQweUFfENt5J8a+WTlec4RsFnhWazE9XzzlupjQ+RNfp
GiHJbH+jsuGaTCcaVdNP1hKan4ywQ2Yu2NktmFkG7hGO847HzK15Tf/buRqoBXBb
TrwfWLsthie5rVpCQow/B//0iQFZDAu4pQICI05itUqU+6x6xzWLbPf2z20cjdPp
eF/NikfMN4qD9i2zOixtsxtzWUe0ySRhkdyXC2Lu5DWUTRsKwE7M/wUUbnHgCDW7
Grk3i8DFVLxaGnxrG+CsvAuEXlVEjqitE2wo8JGa7yVHqI6lOIm1+seYWyWLTinR
9fROEkgIIfzSlCLeHJLXtgPkLJJhIdk4JahVNoumgg9yI1G3lHKg7Y3ec3N/HuRR
HeO/ZMES51o3UnnCObmiSIhKvZe9h0EafpsbBdody8Dvx34r+2hJSdDUtZ8MiYST
HKEoxK7sR18oss64IpWjIactAVBujdYEg1rzWFf6fHQ1z01m0shfRnKLfS1ZGrKM
HQ4Z0z6//YfgAC7FAqCop/M/kM2/UVNTNX7//IP6nsWlA1sIlJUSMxRKE8IrRSS6
CSM3uwu05P1Ags4pgk2tF8q8E/3y8Cy0LhJ/iQJPedooX+YZhvsH+uBE9NaUuWG1
2uQPd8Ho/ZlseU3RjArutX8dbJMpJIKGspbhF6Hy/puyv99Apjw8WJOBWIl1g21b
IraSzin8jUuiOG2tWBTZ+Fa8YwHLZFEcDsTFKEdOROqGg2pmt8q+33Yu/B5/DTHZ
s5fMpxwcbk+oknfdRXUh6ebxkXsxsxwmQ6JozPAdpjsq2C3YUdbLbAS+diGABbg2
T23HKiM3kvAZ7WJm+JqAm5rAgxlrcQ7257DCngOwjkJhR8fkwXIdPTbbc36niJzZ
T3NWtuGc5/KpoLNDRp68vEn7QGDLS6Qbrx8wEendc3X2f42xZM3ZCYiBvR7ru9tW
mRmT6dJ5ie/cXyi3nQFzKB7dWtdJjp/0qdy2XpjKVGP5bENWW2NBHIO3TsskC6my
HW45KGV8kLZ9df/U8ssh/hvReZ2uXFMhI6Ys30Y70nN85BHTog4V1i8jDPiO5BC3
PTIFckxBw7biODSUxxD9iq49AJsuCzYQqvP6+q7joC6Q2efLRvkNI4X0V6RXCaQO
g/qjollvuqwHfPVNeRZ5yfe/OKrHHtbVEqGez41pURuiK0DtVL35LslZ+9GQS25f
1SigxVTvaxMykeDg5mPOcdfeRNJzje7cRLS6WvQhZ8j9EwSirRETixJTU7w4O1Ge
qLENYHKkGv7UQJbdJEbhjtF7HWLwrMU1CEjA/W216bv6C1LfH3mUm4VK//4z5vcr
fMSUiJUEF7F4J6JjX7TTaBjLdiwMBGakzcDAgk5z1l/+Gcwb79yWRYkxkiSNtitc
RGpdwA9iDCEH4MuUJnDjxaQzK3I2iMvjPRxaVzfifYHal1kYMrZLS402lrNQLKsV
rYDwdzE1gt7Wn39c0n96JySL5Hgcj5H6GiQ+wnX8SWMCDrgl+r+JMrXzG9x3qOf3
EOWhZK3Jil/0PnYwlU6fPiE2ZxpsWbLg7gb8S6emBguZYpQuMiRmvuTvTThJq6Z+
hhtycSgO9TpsBGRvs12b3nzpMHp5yIWLO8AYqwJxGBsTsKsRarNuEq3rnEDHRvJ/
Y9kL+PIkn+/4MyCAH4lkRJaq7MG3KArj8ZLp1KSXeVS1YoxT3PYQvcsjeeRnxuVN
s9YaDxnLComGIgzxlnGN+D96KXe1CaJvuxMBe88wf+uA8Y8JeOShBOJAI2pQZpel
kE2HKVE8txUuAbsHZCCaFsWR1y4+nB3oJtWVsDyI3Cuihj+BjP4MceEFXiNtWGQA
9v9gTfQkGeFzVJ5HPNaR+KilErdYSDaHZgoZvOjUwP52gZIT9LRvXCM0fxh71csD
CRtDKKpLjbrFJ1NlGLvIg/4pq9XEhwWrkhvQ/xgGdF+S3B+HjEMNPLf3v/V8dPk9
C9ETO4lduj+C0GdTx6Ojw06LeURESifwPLF0MHc5njSrz2V2fSL5udWUgnurSFtL
o87TQxTao2s0hc7QJIc2U2+UeVRLHFtzWLWxFxk03jyNrNahvCvcg1yxpoYvbux4
pFPuDMWvn7OVy1TJw+Q5xGdSTOLtDxuKelP39bIvRGRemYPzKBJe+tIykOGvz7yW
h5nC/dwAE17VtDQVcRUb477upE4kJKvGf9DU3G9Vq9s+/DifIX3mHY8efIigCctX
XPXjlHWyDuw8IpxuZPj6j5gTHDFnlgCaylgsGdtgrwITd3u9+XB78oPPit0/bFo+
4P0hxu7bfOo0iIoAusjsnStGEUhNYJHQRlOkfUXzL/s1XXCyNMGn2uH/pnc5iKRP
9T+mh8xfMM4tHr/meMoerPUHLVX1njQspGTPkbwGZAlT1EfZ6m436eAyKpxjYmZY
d82Xy6tmy+yOHpoLn0Fb6G3WZutLjFmRu2XX/KJSDbl1fzbVFPRs3sx0S0rf62UA
kvwzUZAzCMp4NsaxrxNn/BfU5fwOV0Q6v2Ytk9z3/kqmhu+YxmXG0JUTke1d6Ee3
fvW3cuHKKGzmOaIXDgEeUIed5OfN4sCxY55hVE6Rm2dj3VPf/edS6rRVlP1ssyqV
LHrbeQ/tmNyqWGAZpTJubVKMgk2s4sbk58QsheHtv2oJIiicVm5Vpm4QhqfrxN/Z
fd961ikUf4PMjIiCpsj4++yuIvl4hdS90E8lFvb/UVXOa9hUlq/sFw/jc+hxmAru
0ROcGIAI0GMaldIW8RVV5vzeoOW69YVTsCknZf0so1512RUZMTMOAsf9kSI8JRoH
cG1qN0/kNeOt72vhGzhZG+FYPATxZksP/H2fvVhZ/IvxJ2ZMq7eaxUsUrtCPRc6k
SJErLbuKZSJInzN86GqZk4xq+viMquoifJfEvmsr2dFgJ0dJ1UDEViVkKA+QyLsm
sQ8DxpfSfzhXWwDsHVgBcipInDFgGKD4JaGPP0+RQUJj8aBf5QqaK5JNG8tEvFdl
dliH+ctugEX1NO7nkXwJLnMhnGTtx7t4TVrFLuCjaVnnc0q6WVx/unuYdeXbnu4Z
9zKXw9d8qHJSc8GhOGZLr0a7pJqdwSCKolnHjdI75zKvCOlyRTuI8VeinBlFJUVo
iVFeGTuZXHf3WAi29a2hIKBDQFXs/+TaDkKSrmZjeGDcYvOV0kBQze7GowLBsVhH
N6oLECZl8XMOqU9NjHb6TR2scO8PbYaYs7LzHRWfOoHGmtOoKX6s8uHV0JUHEMmU
Ail3Cw29CKPXDvVl5jIourLElvGDTKTz5OLP8QHp2nvp1ogRomPx6iTJrlFCKRGT
kVEkj4ijCL5yq88Tjn2PyzZJ8+7uXVZqHRjHe0E47nPK4w5Sq4VGZv2VloC+9ga/
jB493pFJ4J0HZeYMjWaWU502J03QjXbJf5tY8pEe3RaXin6v+SBs0kTCE9ilx3Ry
70N6u8Wx/zFGxiXeJ9sFjiIKEqm1Zx4ymDKmZigBKDrc85oZd8gsmqJLSEw7SvW/
1AW++NSjmFP/liXET169qxvpHoPrFGfBGjaRzuvNWQqCLyVekG80kdb9OVmE+t2s
rnD3RmdYtiI9cU4akYcZ5+CLQNIIjX4Y8Wa94hEQTrVsgk7EARI0Sagvc8S0VsiQ
lDzABD8O0xvpQck3vnB3A5QM78VP+eZujuHT9dZbahfX3rKQOWehGwiIK2lu+itt
NX1qellD3Q3ouJEy1i4s3GVjf171uX2ChJAZ3a2ZJy1XAGjYUcKfeb8aS5b7Gdru
yC1sQbzavybA0CUztWs0ytIP6vxzw9CXeQZe/PnpxRgN7c6fVRpydQ4ROvgcVC/2
E3SnRFxQI90hRUY6RGIeqLOprt88F/drbsF/BjDWv3VZj1AC7W0znB8e1Mq+Ztcc
9RFAQ5g3HS3IQhHM72ZDSPGLXGSWjB/wa9eCaKMUhnCJ5L/mLiZSZOvfTtsDjZBP
o0JkeQPEkNmwUUrrYGXUVEbqXLaG2a1qFvAvuhardGhD/NKqEPIRh7Ey7P3GKcF8
stMARKf1lXckCbF7ibDOlwvbNoNZVFXuhxUdu/CMVNsGk9DgV5J7wm04OZ7eYyj+
CbI3lGPI6K/vYw3gW3rb51ndZsfl/QAn0j5A569kscSRJTIAJi9Fy42Gl8vX41aq
NuMCjvS3K22o/XwJ8VtDba/jjVr/36j6naEo5GdFo+Izv85iDVx06WfGN2h8q7yN
eySy/m94zdus8tXIqAKg0jQTaaPMXMsVHnERYdUPutOyyFl6umfqxu397fswTmCP
ylvvFIoiDnYhzjpkJEt6IAAhi1YZDFrvuw0K0PaQLqqyn5RzzLJ5TM0Qz0jyrpiC
CVIKucN+mHV1Ie3S9pNVQYCTaPlHmd7pI262EoTuP77DJNCxMaQDBXb8HmJkh6bv
xXFs3NooMw+A76U+wL6x+jualmJxZskgfQ4CKx27mmAAuUY5GfAfX4f5kJSRkfIQ
UIytgPnqqcMiVRWEPd5jHhNLIW+YCty2U8pnm0oMylsTBGjppblNYHKDnEs36ChP
kWaKBn98COvmL41VLqv1iql/VmBQCptjQDCfP4LOtnwbu5yaiICiPFpEG91FSJdt
Ad/DNQZSmrTb4mrFnEJsdAsQ2x8nOuI2oNoxABDy6TDiLBa35weatpBduwxaAXKT
yNnDESHlGVILXdPTrRg2O16c5Uc5sXuMcGPfDBla9FuFc4RD32EDR2BdULMmebUc
VXBP6XQU39ManA6e5agx8RWNQ3+yIjjzqKGRKdPFoboZ//tfatGvNmarCf8fbkcy
56mjCOCdLS3J4sft9VJfo1OGbSLdOvRqCDuQ3n2twQ38wNxfpSYhSVlP2IG5mo/T
sLlW4k6BmsB2JmUvMLtw5XTSa9WBloQ6CXV+wABvzI0jGZNx3uLIDuDgCXYq1lgp
i5Qi8tZ09WDHDApxjn8kYnmPYqDQQtPf/3wU+YyZeRqNarfRbjKf6sqm6rlMzr+n
xD3KCLpuRuQmcp7PB6WJ3WXe13Ff7LCjptvwdw2aCbwcAzflNv3xaGA3+slCnC0E
GCOA46QRlMs/j2mlGhP0oMPuEyql0VhWn7QVWs7Fo+fFp7QV2y9OcZhzbxUOiRFZ
mMCizdNn0f3Cann0ax5syv2/JILxyTySzzikqHnLt2fQqHqw6PMttBXUJAlZYG+B
GZEGNXVbEmZoiZBRzd7CvgzaZxRwz7pexgUQ5xRmRElqmBtQciS2tZxTgQPh9OeC
mYDX2cHdNjCb+RwCPEn6khUCxSBqIwB8Te6/AGJ5IR3Fq3tFGnOk8kHAIqseQZOE
JWdE8AqdrXjwlzxStgAAfpv4IZKxJEV9mkTar1+/P46hYVVJb8armLvtnVC0H2N5
5G066o9pBOoo+sas2KZrZo2GBG1/qf3UDZ6XZDC+T6ZjuPEFF4NZmBTdk7aO9h3C
sca1l8RjWAL7zJH58kyvMp0n9dCbgGF4aTv+QPRdWMuUSrY61vYTPe0S1jGdFTId
URtoYJUJaeTk8C9a5jkVbGDlVcAmnhxwRGrGogGP35I6wAiD28h6Orbkg154bzC4
iirNeRk2zzDvRpFyErg6ibj5DjQHoUU/8GaVlhTqI+B6nF8+LM1Fq3T/MC4OJoCk
JWvUAbHaX69weTY8y2hRCpNrir5IPuKC7W2ER3YJ8fbSEjWcotC6z6xunWkUlzIE
ELeE4lKy05BLVucMDrfFqYvExHQKC5JLxYa8Ok8QMSgxeVGY9xeb2UmFkS76oIPt
q711qho5s7NfQP3sto0olGr45duGrBIBAvDARos3oyFWeakoQ31YN7YzJv+FcEZA
sewDp2Jp2X53D6qY9Hm7oXglPMCsg+TmcWlvVdmfUpl83S+G1KG5GVC+chNSXP4J
R/cVKF81CRKp6gXrqan19HOyUk/0i8RY3Ilyve8wRUOMq5jfOa5WJCWA7AoKCH5p
qAcpahjhla2cMrWas2uq3flL2TsJXBC44OZKCnQtG3Ni8eI/OCqK4vvrL8bx6GpN
v2Cxre1wWLn/l/6Tjs/qO6v+cBqgfJIacuy/vVdzJSu256AIUG7mEv562H2BzABw
KwZN2zmz84QggyyhETwbg2rpajMr9N5lcLbMbCSqiNYSzBNLIRZjVkb7X6gi/O5H
7WCjlnW9Ch9CIH6IQkSAtlALQKS5aV3b40Z6ZXMT+JXh1nEYVXZg7zykVwyy3KsQ
PVQhMyzvI9/5VGH+S27bmEHNIIp9LENZREe4WWFC2vKiUszUyeVnhzvPo9LFldaZ
BPh+pIeZFpXb/l8csW3x5howCpViIA1EWgiXWZ3zzB0V0dBIbIu4T3lEgaaHYUy/
WH3i53NEu8D4q2A9lAjkLej/W+FIA8OLS9nZob5Nj0CD94WyOxBc4m6yqye0MVW5
l2Rew1feF9yW1kyTNT3RuTLE2Leituc1RuHjsBdX4vkUXvLF8Iv2OrndH+DdY5Nf
b32ZeLYspSFssz1Q3bb89U3EKd4EYKQBsfS70VLeHSSz3YF/W6tQd37u89xKfpcN
wWFWiXeaxSZ08pkKgmOx9kwwZM9D2AlWd//xKKKX4JV2vZPb9rJZEljb8whdvYJL
39rFR37HnipJc24K/lcNXl+RDxg/3GTfqMomfgHYXxZ3KM9fyUTdwXGjpmOLgReY
GsVIPKanDZ5xfAJ0vyRNOWYa+38JWKoLYuoZ60BI9VibEmw0xLJlSApFweW28AuG
hDg+Zc0MS386GdVHfaggSkFlkCW+j3q+JgnQzpsBrohfHWOj+BHlDHnYMBel5Rhs
5j8znNdECHYJFY9V5jmel6oatA0agyeJ67ertdqc08WLbn9zVXyBKNjklAnJ1wSy
P+9uYmzz1W2gb7kNr6Y86uGxNQpFpGa2tHNgVYQHDN22OkKciWUyRNV3hAC7dMc4
aoW+uTpyh/hfc+XWtstYQ+01wg0XKc8ahdKJq19vqKxVRpd+FQdWQtZybTy++gu2
0n2Mja9J21UuH3zuoMxAnSH/FnmTg+aCEGz8JnvUi5uRqaiNa0Z4wc6bnH0JmTOG
8ZbLT8XHKdfK0Fr5L5RPPcwc3hPN+hwsbTsCyNuzPb1MNXYT5knYzp2qBXBi2E+8
hgt8Uh1dKcdjfqF7sPqB9ZY2jF6gh+4ShQyxDUHSAXBgxwQPAFmezrV+qV5maA5G
99bnrX5/7i63jFtGsHBUSGvayTHVg8oJcTz8dAXHaQ6PhX3GrTBJkuGOZQCHrJIf
X2Y8y9DM3nKX51qmXIAa4emDRarBqKDBEGfZ2LE78YR2qAIWYgaN0QQhKd6nIEj+
FxL9JTmGGNKq6g481XgANsCkc2/LUQUaIo/G9PmW46WGIhifpYCjxwyE+lejIIab
eUxbwMLbuN50nJDS4veNeadYsyysPYlNNVwhhq4Q0Ph/BywWtQ13GxLtY/0/8z1e
uiMoW/nBtGgnnXGZLYGnVE2l+q+AercePVRqgZpLHVJLmOy0mFe7QStz8lcu5THn
CNKBNCHSc6WizLshmI3nqeQmLLjEy2JYA65AjMOgKZKEzHAGFi+j1wRdsOpDVS/R
bJrLy5H173Q6qL/9nLXJHfsUd/SwT6+cG5Ss0Ho3+1SCPuV35AucEr1qTtEWirFz
m43inx+svYdUK7aeU6s8Gx/v85XDjlMNk4QYaj5CbczzRV+xhoR7bU6K+41/3TyK
T3SupdEjbd630UoxJkiWy0t5g7VA82+63x8eKCWM7r8wHyVOUVkOu1lT95rHYHUq
vjR/tnJ2/gDoyaGunTjD5Vp24pk301L41PydF67aigrhq4OV8nZPwN2k3Rv3D04q
bBEKQHM+mnYo8xx7gnuB+hDnT9jPI08JDLJS0heinkV9z741N/EzsfYWf3K8Tg1U
GypUrBukiIH3jdhTsEQ+qn/rvE8vbQaO7p/OjgsnJsgi1chOwi1HM0zA49rqxdbd
xN8ath/WL/3vrz0kU1Fqd4v62S/vi3ev7BtPxr2bh6LVB01OC4j3/LaoOi+7pJ7H
9NIQUbDodIRBAOveINEpw2WRx9epS7sfZAwfPxzK7wMkEd8E6wIxpSoCVxQ7bjRM
QAbUvMpy5sS19XlGq57tIGNyJECwVNsmZNYitaO/2nDiJY7aq9CbVL5x1MMWPPC9
9YVPQDlMwftuPucyrCcKvNq1NpTpHP9mm/KrY+FurH+lyXgFV/N5mNfWxY+01ZYD
vQfxp2twtuo09kuHaoFL0lL5gq5UOplwNz1kdODxHNneCqZmBhTxVKLZv1nv3Uac
1uOGVuF4aI4scfyNn8DLy59+zH2Nu8VxJR1m4z5amb2fwPDbkISV42O0BOYxgNf2
Lgj8wsISEK6emLcYJ7q1CzZUQUjxkTNW1Kbp4pQTnF6y5jE+icDw87k9UASzfbwu
ER5ZfwIM6ESog1KWf/7WIFzPbV0fvrdsjs7fkqRsi4howF2LNMk51v/BEaQ5/Aee
q6LTdl7av72eBIeAGKJLiyZqRoYZXa/iBI8LwOcO0GrX5ZPxlzSutZmzJZgWETz2
UPV+YF3PM1mKsPub6tSDKxjVmg31RVMXA7Axfy0KRYj5LhYiBT7Vq7HUoTMjhkmE
ReIQv5yVHR354CT81pFgT+NqB2CGcljYgjOT0ZrYuke0LNJ4Tf8FZruVVUPD9iZj
EzQFrWf11zWoCXatE0IxbkGbFNv/qGOdw4bChWvJOngJCeEAAqfFxnlIA78liS6w
FwBFERQT1g4xXUtgNOAWHFHFQEmaFdYWW2FQcQR5YBjbiI+i3fmDowXpp14G7+L8
PJ44wWKmBLCuJ/x78Cb6PaosjOo4VDLXhwYdCqiZlsECFksfj3cB7OG/OEAQnIGM
MXvfNt4/WcWIkqMnwtuVbysUqf1apx+piEnCFg1Gyb/JORGPY8lscnUzlV9YDDn4
+bmRmxt+a8Org83K/pCmUyZ3eyW5VprUdN8xsrsbpVDWxVa2vQvNHZQ6b4OHPR+l
9kjIVRaU4e3iB61tuvOUhcCIRX8ikvO2kAc9/0fSR5R5XTX5ABc9iyDxGNMaE2y2
IlV6ENyLKh4R0dYZMC8Yz6QbzIb0KdgkWEAl2uZKPOaDGJlTiL/EfszpbVY2Ceg4
1HadYByKYU3fOUJVh3uvNZznUHyQf0gIAUQvhs8bB5TbdRCrguwjuAgNWhUqXKAP
zZp1EqbkKiQ+1CSTdEvqsUwu50aYf9NbBdvBZu4EtHodj6oqtyaAAdvS41NxYcMr
dDnfgLBcHGnpPVG6rIP1y3t0rVSarpaLECCCb6NmXfJFljnMyG1YtAeS2Hs8+XNg
Sil7d6XXlNl2AY170ygb5T8d9d7d9EGtrQi1uTpT76KxBBoefzfwxQ2kgq6gs2Wv
qUoFgFUzfIhUT1ALP91o6EIC7VPyLv/wEqbBvAw5wv3JfTZolhcB3v474F9yGqJk
j4bMLK+8q+ojkna12cI2DO0VjjACwFL5ttD+Z33+rJe0zqyOicCQ1NVW3RAT9NUp
Xz8Z/oNncul2SKxgq2m12YyQ7ZqZ1qOsB6tHIy1UsWLNkVBFyGz62LkLS5zam75+
A5ThI8ki6i3Bnt+ybpsm+jK6ByymVBIgHMKOAlDabgEj6rnvQvuXT26stZYYASdF
ymRWxXUb6RW7IKpR2JXmauSv4eIgjAOIsqdnpleNj29eXdQT+kMfxM0SotF42XST
lWWxMSS6gvawgAHr9286oWA9zG5cgwTtwSoiyM2kn6QYFjiMHk47OnAW13YArnyE
jmx6h84aIz5J36pQax4QWXShhRCVRI1O6RwgwcSnsBtFRI/zNbCFuXKF40OHFEsp
fNMD5VI1hMKE6snZeNpDQz7kdzNFRD4Os1NCD6A04Wbh7s5gIFKj/B4N4dNbsSxy
AHraFPM+10qrxoxm1IGiI4gxx5tKP26gi2oQSJh3X5B7Mxc/BHpmot1P2QY/hph0
d+Z1DMPlCryBU4Sw/cNZzsivbsfTuZS08o/av0qHeS9qN8LLMOVkyizMZAREMX9g
fr4+/RT1mwOmxxiVhxfCz8AQg+JOlCyndKHyfxDYolF7Hi/GJDUmm+ZrKofmlzgO
1Lw1V8QO/5Xy7VtpoWFcHfiSBfwsabz/WMTOHy4HeusVzXPaF2Dsk1zQhnRaZ2YN
7OnIYQpP8AbaKcJOXk+q3eIRnGR4Oeh/TtbK/CZbYcOP9cjonUPj8RY0WJcrmU9o
5fVzWFiVJiOgW+JOsqSjcYmbKr2u6Bffol00haTyCyfdvarxqOTTSavPMGzStmhq
CSXzi2oFtmIy4eJbj1Xwv37auGUcNgkMB6KvyY9tfTm5siF0yRtuwDLZiFq5e2vy
yUU/0qtP25KXjaWs3SZDE9Y7v+IorX5v6AdvKnLM+o7O7b1b5+Fxp1Qb1MDOeSX6
DrZfmoSxLLxxNQAJgfMXI+HfGjSPg0G6IIuokD+8u+6ngJWsvk0agsEVJGsHHFnk
vw6Sc8a6tq6p4q6oXZaJkB4IEz8F62L6lUgkmeVpjYHFpZTn9LcquFTti98boywb
+N9FcO7MO5H7Na9lSRBR96X4iOyrVJMA4FbpSVC+NCrgeRM1YCB4Roe0JpycDhi/
7XHxw1w9EhWj4UxU587ypg1vSnjctAffQyJmpmpkFgQLkwmJtxZ+NHU++pVgmzWj
J1+69u+2yNjpnNA6u1oWufNi2GBurtTps6zoSittKhv+RRumsx9gqdR/H8x6CYA0
u57031Rt3gFj/LSQsyHbJnXrW0GwH6n8H9CLIjDbbC+wG7BpBFj+CLeDL8bIh9kw
7yYICTkohK3hwK0wsgsyBkiI4FjTAYm0l9bQWK2uPA4Oby+0zMH+rrNeGOA7I22e
PjFbmbFL0FcMnLe42l4QjOIxJkS6n2vLcYVSPJsnqrOg22c9vxogA/j9rTB8ybQW
uENbh0GiaSnVYOKTkzqtBYi/vITcXcFFfHnZziXw6PEDb8FzXwsskTqh7usmw5Ys
nIXZkjX0ovsHdcwRPPHwOUusF70nsZu8O+qAq3xdpVs8ebzAs8q62WggMD5yB6v7
ZoLrJEE6yCyIrL+0WAugB3BG3GBoEBzRILgdmtNXkBdGM2EVfWBJs8ll35qqHDgK
yzkykdP4u6QEgGhn+2DtrcrCM5O/PQX5nGx58uOX7NlV9d5gUfGJXNdxHezQYVjm
H1qHGr8k3kDCZrgb9aoSdqy9oF5jceuGvF9Pj//ux+5tGnPd+py+LmvYq4Ak2io+
l+waGyQkrMG9EUAdPte9EbMT3QoEEWj/0x4Z7AKOEmWr+PclBUiBAurohdPJZZTL
VOdyA9lng3PJtR+bY03cjWlyBHyi8BSPW35P7qSzkgKH12ezamDhl9LjuQ9zwYCj
MthQsF64VSYKzyp+F6vKpSHqVd09tS+tl5YrF56RyWm4680kwASz1pkZhjs/IIoo
QNviHXHWiRJgqgFDl0eaYZC5Zax/NtQ3xz+wBx6rQVSNv4IGIqdTq4cw65OQtkSm
027LmAILRYCkcFFioxhiBKcP79WlyYvLOMlHOkfMHBAqzFi+hf0UPTOOMbEz/WnX
ebStxaxO/6xlv5XAjGdvG9fYD7mdWecIJPlEn8yQXOmOScB0H8x60B3Kud++OYHr
2acD9qrM9sajCDhMiPagB3N9D6/C+tM63sny30SWw9ZALr565iKOY1J8jwvNzATK
JL0CS/iylZvS7monHbnqlt1S+cEE0MyAXL87breYQuBB8Fgtjda3ZEsu5raOKu5Q
Hdkt3H9oYjZbffNiulRnVB41dfI1jT8nDNz/DRV9dHgkw9TKDFWZGa7HeXmVMnzx
+B1X6yRfEOMiSQagRMGL/9YHZatQGWCj1m2DWuCNTjBrCtqCD2sNKf8BhjP5EHTG
DXLGiBaVvDAyPCeHPAJyt6iwxUkofO+YPwYXLwWH03XHWtK0Ps+uw+UQEj5IPi45
dhv+bmnO4qz6f90zJeyDHBO/mO0x43zRRbOygXA7I1n0g9xhpTw2XHGut1T0Oa+J
S5EBbT+UP11P/90kBbkMW4zRZ8nb82LZOpHATAQEtj2lmQt1LlezSDpcat/hhkaG
dNo/mkgcxfhkEgeu+rfWjESxKOkB1SK+34OOrhOhHEm223wie2b/7RDwwfudDxxv
olxRXzu7/dyDDQIgLPSzFiOkF+T+ieyMwjdzza5g214GnuCvH4aCgDtvWAUytJBK
bIjYOzvqOCoT521SB5q/eXMqejQ+07aQnG9OaTOBGWj0o2a3juOdsVjK3MlVmtEb
e/jId7u5rch6vLInOSzQgJtlW5EZuTLQhi8DMW5tZ17zIs+9YV6nFqL/o0Q3VGpu
vyeOrdt0qBDxTgQyHkCsrHmbW4rIkUVnmw1H5Rsr4/Jq2n+DT69znMEJshgY4UdB
dKA7F+hmWXvcPAtgQKQKSlqc1+Z56QKy7n8iDoheUyu0g2vhdrKPDAtx0ecdk5Ov
KQEn7boHTQfJS7hipCAUXVlOwv4L1QSEVkD2Ea93R4Yjbr80uvafSEJ+vISwJraR
hiGuDm4lDxfAu1SS5OEmvAgnD6/9bK28JbRjKH5CKHNKUjMWKiXy8CqXsTPEycCT
QLH1PDAIaxCeBzsz8FpUJKh1SVMwQHLWizggx73z7oThaBs5Y8+yXxaF95yA4RG1
/5ok6/0EbuMjL6WWBfKdWQv6EUlIeN2ho6xlzs940++1h/OV3w3tQ0GSb5+M01XV
a2KJlZzn63f2RpUNaLV0wZsvQKyYOGyD162KOZinGBB4ART5Yvd/vPAEv9Hjji8G
slFwHSFOOOptpgN9DFolOtMXAJz+yyWXYzrbjxVe80yDyrzivIlo/y32Q7AS25w5
Rkj1c0S/veOrSG9M6iNmQR/Mz+5whzrl50nElQTayKt/ajQuhtQ5CMslQ3v/8YKS
R2qlaawQ6xi0wjj7HdrfxP4OIF++1A5QcPqf3LjXENPLYmts8V7WbIOIaruZ7ATR
yBDk59hfFICR48BvsnTkJPSe1jdYRrolmFyt01+6BJCrENbXo7uDaooLIKbdhpKx
LiF6A8PyQHOy5P7xb0+ddgcGPCYKVV8gfijgLFhZcoo0kmhSdd2+vB56Ravlvzq1
FRtw4d9IbfumFjkYxO4bT6iEVELLO38yiwJnOCUqWe1RNMqSmENoQpfsl2/WwToT
GvyLW7CBMDYIAQWqOYqXS016qDzOWzCwy//fY/URI+RkNEaMx1XLXNEndKmQ7poN
86QrhVS0iQ9QUfM7yodHGy50qvzX6nfdGR0RbaYHjDRXMkd0nomfurjA8saBYHLU
QqM9xu+CjZie24mdfdIKmQvfeeHf419zktlu5FzYs1bWMoVXmdRjM/vcurOFcb5d
4P5g/wt2uwjGeX52ZFUBpeqHXglvC/VJ6pHiHHSI/agfUf19n2VAi+cRycDAmXL1
W0eSYkMBH5hZFe8+NCiqL7VPMqSyox18ed808v4uUyG5PblOhITZyN4pzi5fzvmx
XdiAS1kG8IMe3G3wPmXnT27O9swP1RnC3BkuJ+SiHbJ36q4A1+DgFgJ2WgqiSTkW
ZHLBdKYWSS3+XlkH4MCu8ZXosW00AqxXBglP8BxUKGiXy5SWjfHBKLp4UfvOnl8J
JMTPa4KX9Nmfg9eZeU8h/vLYw7p5PQAC50FgwLrvnbLbT77di6piq0GaGxGWCXaC
6Y8FRVXEQVL2bnEtQG3PD4kwGvhJSpihwEqDCCvtUrVrF+fHPFDD8anA6XSrPEOh
9XtiFfJvdT/d2H0VJvE1NeY0M62dSc3VSaVev3Ckln9HBstrIssp6MA9jlmNO9/3
/SC8kY7aV3pK9hEDHtu5AiFuehHhrrf/wuB9J41RsznQ/rh60HLAzjBMCzA7Tw+H
w615cIffhh46uTlKv+CVPuTrNRgjA6eG5+jnUU+HkrwHSOkjU/wak4B1eXoHDu1A
RgWhR+UfyXXd/nGQzULYi6vsaag6pmu+hn3Wr0sY2H3Ga1xqH4kER78pQoaEUhsY
onRK5Brlg4tjVmq4SDXUw7zE26/13nfmty8nwrkfNQ4+ZhxFamPOEdRC2U8RE7Os
JEe93zg42/waa+pPqZP03uqhz5102dXGyGV3IBwPCXDpYassWioWIjWyMkGOcV5z
NdJYSITBViPb29ddRvyTU1pUNEqJImbT0U9c1CDapjQ3ryWZyosXDK8CcXlBnsWA
YK5Joj8anpUTBymnRSZ08fSoA/eTPRbNgxQZwGQI53aJ5Fwud1l/eyXlRt+6jJrW
Mi/eeZmPiqWXEHYBWS/+0ZpRpzn9imqxYY4cgL0JbqjsDC6Ftt5PI0+GDymssZDD
MlTcFmIS86Vx0euRA+GIb4+G5LSuvS3xI87uYzlgIrUc2zBkLCGMemA+RMDYi69U
B+bRkAYD8ai5oClI2NACLBYPiMxeAqKxSQ3fhiVqh46J0RcKsmMaqV5/OykLVsAp
DrLcrj9fozn38/nAJwSIyO4BrZZ7Ox3M6QIqdLzGQD60TKVLTfQQ5mGIEf+kGv5E
XB73pDfou1Q3rFR15mCqUKOSQrWhhR4rtRvjvk0PFc8hGU+pNB7XS7Bu7TqkwY99
Z+JDhjiB4cw0zST5PatYSLPsxKn8IFXM6EjgE1YkKk23MghWFXLtP89QbJcYVshP
AoRpg07JR6VtjJT698SHAc8Bpfjj3oYCHeyqazwkIRVtD8DD5No0VMTZzgJG2X60
YAQhpaAyIS7BrlZ4bMeI9eoZg3f1pOsZNzajZQlA800LS0hvzjrzpYndHi1lt4n7
0yKO248qqywNK/IznCzPRcoosheKfxWUKydXuvIFPRIZKhetIZpiGUblaAqf4ot6
DnqXUflajHQ5REDMXpSGB/05EdByHm6eZrLoJow+jFZ1H3s9d8Urp9A9eOar0OpJ
XEsIt9hqpEoM3jb8MMn6SfQFI7XmWx8TZFi8tXg+auE8k2PcpO47xhEo/4PqUIo1
93RizUUlpTvaxh0xE6Ek2s2c2vtDeHPjhWSCqrTnTAlBiYlh6pHiNQ0bKzU3ZG7i
MaWvq/lC/+crsH2iOOy0Ti/vBOMxnvZcia4OevB2cdrvaFvNykqIGVq17YKHacke
rtSx+iXO1r3bfueLuhfSQ4eE9vR/XdjUchsLl/z/RU4LxYZZHvss566nkLNRhJ8r
aHAzRJDbf81WascIAO5ZEAIz2FJUNFFLAxFc8aZ3bXsfwVE7q8EvlatMQiPM/yG/
vRpP4MuoavJko5THXByqlO2rKnpMsNHo311NInM/B00ROBf6ny9Pzjc2mcM+tJ/S
q1iOis9qktCgg/2IOujo16yB20qHIlim8M9KP03cxPeStx6JGwt0zBokCONKxFhT
/qqisagV+YZPRnl6DL+b6CCSnmsduNG65dpWzS4/A4S31fE2afyz6z0C2Omtpfvy
U4XEvgFVvNvxhkYTs4pH52WAzeCiBdqVZKJ60yPuP6Mad3jYsS0iuc91W4lCSYZx
W0PYCnkGL0pyp57nYqnKvUM2GzSqUAF6cDdEwv1Pj3mhtNuub9cxQbZAoxgcGA7G
PtXqxTREY6OG9Mwp2cDPQJcFHrAdNhIfZKJ7YWSlND5p1frM1oCulNtcV8bSghs9
a7IUXGzv3IySWIf/8SzzVRfWI9FLyQycWQ5VV1d2werTYW+87s59QOnbn8g0/Q0I
RMszXIS4ElNhPuplhoB65CqyiXeW8NQ2GIN1UGFmeAM41kPzzvGl2I/BMWDvkEGy
l2/Wa7MO0cnmwkOVrVNQZJwbg0G+B8XHXrWz0NAmpP26s2S3Dl5tu68yP8UZBeKK
Xfqdotr5WbozfBGIpjuI0PK0QgfgVtsqePYRZqxvSrLqU3X2jrG4DCtdd9aVA6Aj
FKIXx07dO/YEGpu73Kl3J6YGti9DPWB2iU+vz1dgFTmTsl8YequQoa5jFpgp3vMi
aNV347cWqUPYM9mgqfLqry9La/ux8vEIxKTzYcpS4pPTXYF0TBqCKuC9qNJuiJmi
l/VHyZqPZLTtiMW3Xpz21FGmtBVnE57ImyKY50X0LK9CREZ7HYjOTWm/IUK+/ns6
RIjwwVlUlayf8SE1JtWDDOx+NRO5HhCcOCn2p72cPx1tDKAPv64aC3RjqSP0VjSH
8LH1oTw2BZ6mDf8y03pm0Lm7yfiVv3EzpmMjb1UwZVr7G8lQhU75T7H4gNRrC1Ak
u2QpP8SSoKoMeOVLMGCus7H352qwYGqZRarJsLgdmD9j6MKLgF4PCHdszL/WBpTe
F5lV38y/LTslPyg5Lnh8KK6gtSED3OcOCXU/fj0LnSRRhEnAO8lsUDWFrpxv8J3O
+6sO7Q+0kmsvgv/UJ+NNVrJR2afD0F1NtnlVOaLFZhI4BhBMwXaSZUQxniI3SNtN
UUpSGGgRtsoliM7nDqIgDFMaiTEbycEryEPcsV/Az/OVdg81whxurXPhios7xdCV
1XMwjs1YoaXBKtkXNtDd23N9zk/BhiS3tHh/TLg2tZgPBxtibHDAeJ38CpiFTvys
i7+iROOIXVn4KgzqsyBw4VtAI1VmHA9GM4kpTz7+xZwUobdTXVqblBgmR05PC0f4
nwpmPEqSHelcfYoX8oX0MetzM7GWytJYWzU558+OPV6gBhWrV3yhsMAnzvLQesmK
IWYMgJLS3Ex5HHGt+vXgCL1dQ0GbLnN0OVxWhTLnaasVq+w0Ev8JZGxAibMTylhw
Qfn5tJIt+DVXGxjiKMhZ6paAI3PFOccMq2If5VhhAqoIV1+hxxOb7i1ly1a6dOFN
KsCC/6m/u3fmmq1Jy5iD6r9oGCtsCca4UkI8NJV4Hs9fllZVJKKnIakwm13eIWCR
5LmV/ryT0CYcuTciOS3fqlxNGefzR7WOVLgEX9GpV9HjwsNBlXcBZ5w+Jt4YiqW0
OeUOGdlffWIdbZBKX7LInXMqTagTXS+QRDTWRegxBjDIBN5fpBcwefrx2zBVSOcx
fVDmeF+i4Mz4uIqPbG4g/NvEXatmRxJTNK0uAGtM8dgJsSs6Ptnc9SxczU9Iow7+
IraJA/4VK45qw+cCgYmy8VoxIwpJFvNpZNazElbU6PxM7AX8RAmegGSHfv/NwK2H
KnOGJPBJxD47pN6CtC72UoJg4LX5s4t+8MiLBlv2IRYRMQedmC0RlXBeG1Bw07k8
a593nqORjjlBcQBKct1EZjk43Qv8fSHJmN5wMk2/l6c6Uk+g9FVK26y172WHZiXi
zZFFEMEj2CazaUdz5kerJRmxo1f+rHxOyWJ/2g0OPbEQ9ZZ3hvFTbo9ZSU78UZWR
B4egHOIG2AFjYQP7v5aUz1QkjIL9t55YXi/29BqQsphbXkKZ8Wv8Af0uaErYrhzX
00rs0Tpm/7KUGawqLhgk3wUqZbADcCqsZU4I++iNcDWMf7YuzptI6QfNI4oAehak
tWNkYhKU04WEO84TaV+0HvvoXxL16csD6FisQBWqpAmL5hoNPbmg4Lmjc7FMOo6b
WFAMhGrJRkvrcsdb9kMOHl3sXUXRCxypVMWu7Nx7u05wnmdofb8OiLhs52hUFtS+
GQgWS3OetmJxG7Er2IVKmxs7jct4MdVxIDloC2qlFf5T56LzbcRslFLsq2Y+vt1O
GFFY3KWapo4hXvyhQgASXI4qhT6Kcj9brqSsIc4Hfzxx+RyZb8aW4uxByeACKa26
JCkVactdQ3kDcTQVbSuHiPfXg9c9EMZ8qTzMT2EZnxjdmuiyniWe8dH/zd5v7dG3
g89b4TMPCpYqaLUxTfYqOjrQX+xJ9onRpgU3vAK/wUxGDjhvtqWT24m/5Q9kW777
meHRGnSu3/7SRmLjKaEdTA9r0flqOhgTWRee/Y414K3bKiNw31XuyucEjrr8XP/I
7hFm1Fsx1GrTTEP+EWEVnHm/jgwUzUellyrtIs3xJ2HUH4t09r4M/sCaR4dLKVTD
nUYd+JIYLtrdWVCdwUOPHVdPX7btj9TmKxko1fX0ytCdrgRtSmSJn+k8XMF5PGnM
QXEgQllkKkDXlOKD2jOfZSJhzrd+O0ML0uWa46+eOFo6q/1zZap9yQJNrylNUgVe
zeQTY3Pn+L8PuehXRHGvVIk4pFJ3tlGrSNmZMZBoKyGQF0YXID6AsvQdHTxJTimQ
zQn/mVYg0GURAnmEWjxD4l9Ff6IiyBZ/Fhc5+6YbwPM9qPWrDkqmGQHaKKaWKbz5
YescEfDNlgpRX6kMlhmGwOGzsAkTahNLuPd2gdi70J/Bi9/st0GnJ5BjkTRsnwFd
xW3oOEluENsN8jJRR++7Dpf7q7eodc2bpt2ENeDDWyg6fPVzFnYh4Qe6ALZg/iUz
hJCgXmJftUV84M6QyJLJuuBMCBWP/spJw9fS4WMM+JJhXkfn3mVAmNIpWQGYDADu
naCMvBeNV/GNR0zpmC00tPaCpqGaZj6vZriAfZfRy5cLVe9Q9FHZCJWUOhXSqqaY
POIurhYlp/o+eZVTKMXzLO2VccDjBGXBKspY56PFLPRt9EYR9fGYuToG2wrWDHp0
TAYGx3WvqOgPuD+ahCVlcAyxxeJDURwnpjBcZUCg84fiG0cjI1YGKG7GOmxzsoD6
Ll79kCBY31apdkxdyb3j1qKzQiAngCUJLxeSQT12JDHcQSXHBOiwXRGhooNUSun/
8bmTzOU/tM8d4zDxQGfTRsE0OZjP6dRs7WiLRheBYnRUm8stvgrguCQLWHfIhqie
En54BuQytrNe6nnYZtooscjzWVR/Dg8cTKN7E9TlNcKz8lIExz3ZyalAZlC3uWvS
AKbVLc8LkGGDWRlvLR7wbj4x6lCX1umhi/AKals+0NB9ArjcajNO0qgbWzoAsbwT
5ZYUs+ma0cz31fFp6cnzbvBdMCkBpohpO0xBd7ZpdHHa+R2/4jAz+PidN5p0i7r7
jeRq27V39a95w+Va4M0u5j6Bjz62nQt7cpeVDQzW3KWGPkXPfrAXhe0741WmZyBE
1Za++1NQiO9eDDzgQFEn4sQD1dtKz+3CJkhqj1PNsOwuEmu1tBFMzU4ejB/KaRJN
H5IFuneuV1qnU20InoyczEtQFuAPYe276qoxMasjUUT7QkkvFPDP2Lzj0oJNNouM
pg3IZhZXcUSw1WIWXpky0OM6vZvFMSy+IFT78w4HOC4WWv3VN6I+7dolUfvxoDZt
/p0/TQOtSzr+3PQuxz6Ep8kZ8UanGRHVvHEhsEB6YkG188MmTK4HYWiv60jjXPO/
fGaT8p14974NZuLIFoSIKO6B44L8K7nGnSQCS0mxLepUjKAWpDriiBw4UDlBGnJ2
Lcudsbxs07aseOPQfArRXdZJaNBPvhN54zx6awmTIEvd5t9S0A8+B5OqXlJMlNZZ
w90ML5gc70qlyRIv4+C3rJMImRaAFm+eq4JL/1SZkDnJCeAHc1Q8h5at6BYDT5St
NelExV6nWI9giUjF8LmwCaXAwWnb1KSF7bwGDEyK2e1ZVAXfj8luGOpnUL8WHHYx
j38QOP367mO5x8qZwbc1kQBAZEIr8dhLEgMnCwVvJNmQzruvM+HOJeNySAin+ash
tJWRPiM/YHrF1jH8Ft+u2MBM5iF1v+u8ZApHW5tKrsoR0v2hHtz9kRkeBjPwfHHK
4oKQ53kcZq3CAGRro1mMRBPdSP5tVP4diYj4CQgyV0h53auWjoh5V55ZEfDletBV
BAKHGVDclWhYBMT9DC+80K5x3+Mm6PfHQXTHD1ME7IdnBLsSb9+/1rA2LYJuo+wc
qCtdtSTXmuaPuTfCFM9zlSLEvkxe2gDp8jK+xnOVeKkd+tyGMCWKx5rzaUyEuySo
r5gVeNpC7lkdSpuuk3Bg2d94+v/O4VxQ+uPQL3cMBprs76RMG1cUcocsQfrzlYiW
E+2MzdBvc4eC1DODDe+DyO2ly2PuRS7R6D8ZC2RhkkZmRIrmC9loHRbsF7qL9D6d
euTrg2tkq3kWNFO+Zw701yVK2KoG/TxnVAkysSc/iUPURxNAesNdLMfXOthi+pBJ
3Lp5ZUPZxAGzgz0XXWi1vbFrnKmkF9pSztorHCRaDxOadqbNN96RqjzJ+M/za+Km
jtPzz/krcW5m1nvImTRuDo/VROpP3DxTMBEzuvyY6Yt+loi8CC/n09d+QZQEFBjG
hMrocVSzmcGuLtzL8PIl9HpUvYNMaWorV1YFpzm4oSFfKkovwPDCCdiLxgbNMxeS
0Q76YnkdEfjxrbnuqj9c9QVj/pF7GR3A1et2nW3f/22spYLnJB2ViHINF8aD0iMo
LrOF16wlpzokj+CIwiATWy22BmEOMLxLiUh2hzMEWJx03vsyssY1Nhh+V8dO950P
QwtXrZfYTaeRGoFsfEVnel3btwQPuhn/9uml5T3NdzlP0a2JE44k7zsrjqS7ELRn
srIf+B3yZ/M5mGbJKEdJcToyR27CmoZokYN697ThhiDt0IuUngmMR6Jn4CIPY3tq
1o5OhPbmDpEncs+JCrbpqt9CDNkqJQyjtfYtcYRB8kvXrLhiQhrKSDyaM0HM1Tgr
ZUZcx2WJid3teCz7BQi9+K+OeVkGr7X95rpI6GY5qduaWMO51joHRG1wXfMtnQ3h
phmh48a/d5EatgF2EIIicvTA+RBXqOLE4h0wzYCSLUsoGAsHjUUnJ6PKJe9uH7Hg
xE5KlvFFcYtOrXSBTQHJkuiohfF2JRWjxAV83vpMdvGuAdU0kY5fdLe/aN+Mj9bm
7ekvcVg0QBxkPTkRO+O+/n0X/CGZD5yB7zwcVZo2CuPqwGim5cY5R/L8YMvGU0fP
2OBBuYr8BDjDEnuQTHHIhZ4WRllJOvqzvh1jnaON21IT2lC8LSfuSDZvxVPphIdz
SDUNi+ce3OC8jDgtJ6XKMW8ap+IXkVVzQDGROFzQ1Wz2beIldM8KppWJX3OxQadn
wbBRlZbeQ82RPlJwRlS33e/6keIlgp7SyJ9jmbNi1x5m9/vd+z7vB0IQUY5bkBEr
bBe+gnFmvMMsY2SeJIDLdpxAODFyovlVH33xtBNd+uMB6CcBIuavlqHBWKgnkP9c
u58mBPJy8mHnSBk1RcxsGjD8m/n7qtq9lj0bnIIgXw9v4M1PwYeuIZmIh8Vh8y7v
gIEy2kJyS6Q1tNI6jRun9eCsiL/cVBHrSOt8tfbiSt/n9Ctmf589zi0MMU4kgKlm
am9Tp93JoCAGVYhhoU4GCMxyYpgK5xliQDeoE2zrZ2JA7fTkKhyK1GquFzOAN9B8
pS4TTi6HmmzKm/4vsX8ZBCzlsVCpn1d8OeBCTegRA6Fqp47JabSIqweqDZei5WdY
hZtv0TK1YT+qQ9YRmpmnCqSc5k7JxjaZRGf91yz4/DCHGn1IeUAAYj6qbBq1K1s9
hi1k0yFUkfu0GaJdeN7PV3zCRRftc3xRrL2GLwei7wOyMTFb6NSEb5Bw9euVmAmo
iisZ72llvz0cWO8a2QWZarfRz1jOxmajCHD6t4b0khH+cLqfiBeLaPNzzBAiGW/r
9G08UBJCF+96Dx7ZSsTerMUX+V1+3ndlyHJjDj2Ck3MjX3EvHAjnLlwWWQ8gPk6h
C7cbf2hGezkb0vi5xvgKqOg+2CIZ0zc/C9/xDh6v39CtEmRdR9BJ7tVx5F719SNt
aGdiMw4znmbKtQyQZC6cDQFMLzv7iEcoXOpmxLUp3B4xpZ7TL3xz05cHv7LuWR4x
kBsGPC9fsqnu20A95WglNm4TqqyHrQQRd8DsTWtAdor66eSCNh2NsIb25DaQPWxG
QOzfjn8tC0wcH67NUjuSyaObbKorQVVCsR608Q/m7LR8LOwQQK2uLYMvLBDxrTLr
txpUpsTmqr9WmhFsfJU2bStPNBhM+H2cRn7+UbeAARKXx1tVvcSnLiE1fMCF0/d5
PrF8rQqPTwZxt01ZFKyjwHxkz7RceL+fM2SykcYunbgl+EHT7j34AFxWQq+FbasO
61371XEXeKzCWIU28kgcaQNPp9JinpKVmCvlVnkde0PVla+m8JQygp57Dy7BvyyH
04+iGgsWnJgrFSKdt+fPSxgpP3NGoncbgbqPOLT67r+r8wCWgue9kP/6oyhutIju
b8jy44hkQhQ6FUG6nyQ6Dve38d+oQZB/vwKNYVHoKPhDcA5/lRs84JSXsbdHmh4i
eistgjLC70NPIcSn6tACCrKGSEcwQ1H/3uVDk+1DN13XEOXBWkICamCxoTKqeBC6
0N8Vb9WlLz8QzwYRuqrR1KGx7FRjE2nty8gPev20HtZL65LeD019wU1DfE3JbBNm
sKMWKvW2g+B52ohYaBVu+CDYR99dLdU0yCWDADhRg/D90ciIXUFEzBJHaC2EOyNi
0lZw0XYg2f1oGsrbMRhOFCe6hudmdkN+fmgD7quZEa58gzwTvD4Au+PbhLujI87W
s3QWwVfjNXFHXEEcp50U3V1ThZr0XNKmBBgliY1x7a2qspD/70w2C7H4+kTKAQqR
q8guxGTwciFh1veGoca7nQGMPuLryY6gI2pLoD4Hx7QtvDhiBxALZGrt3wEdrgPv
F5AxUcX7gNdlFifjzQG6d/w2YXhN4zzxCUUipbCU5ZN05ELQXLjYi5vT//jvUVQN
I42d2Uqrzqoczmk/DbRCfWRS7DqIjaiOZhpegXJDiklJGLReAZzVTgCBciKS5vty
NQTAxRhNI64XJpEZGEQAOUoiM6hg8QQeZRYpBIW7PGi6V0om99rlnAPjdG4rW4TO
w23KBUeMy8UgE3aPRrx1995Ol9fmcpPq5Y2qczVZjTPSZZZwmM8s7VmcXl8HIJ8T
q0qc5NT6dZXota/O1njvJN6ncbYWJw5jb2YRB95sVjmprPOpn5gj4uh/L7ZH5aoW
zw4tF2anNL3y6LXKBs8miB3Fl/JkhlirojNqhqkW3FFCdw2QTbKcIYPi/KWCjfgk
5CzDNpBOekILLMLL+Mqg2Dm3zxTgS4jXHb5u/JpTNc30zBcN8cC7sxSM7tMha1Md
f5v9paw+RREpZoJY68XeEXFDeCxSD2MwH/oNTYinQGT6kblK06ANlAe8lbGC18Rm
m2mObsyyKmnda07O+qAgf3Ye+xj2w/eycPW7sd76G0zHp3w7S7SKvFQ4RpaNks7E
qjSbRJ+WFBnzj2M1/Zaxy29LI85d2k5tJXUietcz+aeZwmcQbEbeq3cd7LkO/f5i
AwZDmDDq6xt45dYAMQIaUapj1+u6gvt5ukIkvVGYVgq3v/ZcWR/WYJTGKWwX0ji2
iBh5ARuCT68WW4euLH2DAFkTbnoWaWA6FtFVpKVarTi3XsMbWxInbBi2KVt05Sk2
FsKtWZGpKsyV5WTcUN0690zcmhN2MYslCP7gMgPuxhAaDmcazoXHUV/s5OmEmbYR
I04+yPAuHyL0d3jcjM5uJWUcJbNhWHAie/RH2casG4m0ZKrQX7f+8MDYj2TedQzP
0gCqWf9TaujIdlg2SYYUFUO8YW1ouMmsoM2TzUXy6hAmVDt9THbEk/iu1DpLrusy
s9JSGuJhv84nkDjEonb4w2upESgcVkizy3YHOjdmBAosq3Qrdc0dXVJzsHhRtl9B
dD1bq6dmN0+zysjNBLlRoEpa9gDgyDymHv0sFKrFR8GioiCPqeBGtNPKxlrDBlWO
aBldQNCB+QtQ74dE2eGFr6yxUeVWUf3Yn8VGavJ2p4ZV8UJQHx7QhiwawYYnNRG8
5ifkf4AkmIgf4zQkKQOa68JmFXcJ9Jbjm97zyr1wd/avXlyODd5Gxtdv6Aj/biqt
2EANi/lWzNdmxy6X6DtINl+QQKP7I366mYbdT1cjP+IGhMDf/y56awfUz1qZKX/7
FdL4bB81dIaE7Q+v72aL/O354UcSoUIqD1uGjVpeK+CynKxLsArFGXOS52D8gNcs
ucYwqeLvT22C/D/wmz7bfthAXqP3BYwaBwuhiodAdsAIvHlz3ANXvkLtAVaN0UPx
7rweWuNCq6a4R7zB7+Fnb7o7+q70oGB9l0jiLC24vv9jac28XbBb9R9eMqoKIDtG
mOZrYE42qtO7SpKOVhuyNy81L7XFRyB2HrqX5WtlmHVyRFTEX4zPZ5mL9ptOHqtZ
CJAcS9WvpIvqCW+ljBOW+3ClbORHDJpKSF3JCSuJel+rQfgfD9FvAYfhPP2Y4ZwU
6pCD09BqA4JTFF1PI7UM3UnahDnyYJG/hckTf4YfAMArOIb7OiDGpaRagoO9g8Jt
rNMlioVaY6q3f+PnJhYuvkhCSGFY7V5RktqoVhB6nhAZs/5Bltfjj+0mCFQxYD/j
6QXFmchC1UIXME0xJxNu64zZ0yODVqQG8zz0X1g+PQpYKkoDAh+4507zNi8w3O83
5WyOl7/nvURBiSTw/N45W9BBOUslOEKBBCoMFi6zzW4EQu0z8Gpkk4ZU/Crfy/A/
eupYnyN6LqzqCy8LPoO70zjPg9dqmoDIAKYsoYpHY6Rh8uQgDdK1eFYagxaN8gGg
Ovv41yEJ1TtFdVpTIUcV5WrmVr0zRBSzxMPjFadyS5jtGCCnW0YHYKy108wgIz1X
Vb55bImTOBBN0INbKygkBa+hShxey9hI8siJW4JMEOpDDgF3sPChGm+ieXwiMMuO
L/UvMQbf63ITqF+bZrZJlrXupr8dtWj82V2M4KXxEId+bF6Ehz0/osB2IRUtv4sO
jluS6oCmZwzaV22gEOu5NJrWdf80zQFIpAg46REjNkwyCThytg6wBL2L2TKXzzPu
z+als98ICZrVOeH3eSfucjfQOp+QJZ4e9JJ9pgKQ2eK9LOhwcteOVVllXvgPdINd
zZOwvU3pJw4pv2bWaHHq+X0MyL7cUUfuuVc8oB+iEBrezdAa/oxPZRP+XvQJiDVW
ySVlFD57QHW/tDcqjnRmy9NTD5xUNAGS+Q9C0J/w+8HTV8+me+0KWJKf8EbtEVTW
0Y36sHvzt3/xWmxdgxnrbP3XkDe4JDKL7tUsJIIj+x1hc3+5a8fpLC3YtTE2T8lJ
h0Mi+xfCdNP9RtkJarT9RwKWf9JnCJ6Zi8VhXtetxUKIcR0mTpXRkHTx5pKJKRJh
RNwh2MwLobs8uJi4FHUXyEqccI7DbL4JPTB4MjnHxFTl1REBoTcYaQrQaOkgoYMb
oHJ/Nw382N2BSQX5NGE1fyzysMe451IA2978W15ItZ1UvYapLGCy4maWQwrrrA9a
FxLRYSEcn0Pl33or3Syg0cn+zZ5VQk3yaSQRPvemdwp7EFiovr1GiuML37JtkzFL
V5s7GzymaEyJlYPRhTsc3ZcZflO2fBL/3pwjzhy8RQkdZCRtXEvyWa7WOFRV73pi
kEXOmixiMn3kh6SeKaCoev9R2CV1QPRXBARjZ+OuIZJZQ/ZPFUg3TbiMXjmsKPuE
Zi332aO1ryWRT/tZHUS5h/mlmqb3OQ/PwjZuMwz/hTUnSvXN/PBMx3gRu2gLNfwm
UWhObJXQ6ErFDM8XMYjAzaZ7qqG5OkNWAvd39Vd+dSLYqmXcafOkqDhdAoM1/Qcl
NjNbjh2mxZBorX1NJqV+V7jXPwzYSv2i7CBhwgFOEy0LOGX+mNB6Dbjd3qa2tjPr
Nso+rN1ca/we/Iaq6Ue/k3dLYSC5pQ7UY1OC02HBMt0pxdz0r0XaNP6I4NTkXkxZ
8IVGOLGSmC0uaLvyz27qEtZBtUTu9VJS7YDao7DVVRWmOym7qLYn68amcFUe0OeD
7cdgYYuX0kg6SvomOFHqqafwvjK7Ko1QJ3zWRV1xPyouXB+BcvngkEez4SFOpeXf
XaHa5UF1dIB4BtoFv0c3AoUYw21GKgsdOVS4zYHMageixgBLNxdm+cMbxThyQ0aW
UP9SFMPRZt+8FoaKlAv7XCmCJYH7+PsvAQGXI2g3qIqXid6S+cz54IbSe0eZSn3O
jDkIYtjWgng2zomjzVWEbi4of6a9gI8Hqk0lt8+K3ERljair0lx3cjheOivCOpel
eM/MTzWnMSb4PtyeQrqOU+EaRdqTB3aB6jMJv8Y9GmzBhQXz2lvT9/OZHE21MUcf
Ge1xD0aAbRrA8/FU0eR+FBdFULQMyX55yVxvIuAALy7dx3i8Vle8JLEoKCkK4EVi
vOXrjpNQL+Xf016JowKnIjD+6wKcPvnu1LuLYbSwmBXB+h8KHtmlK5dIgHoPLDvF
Ym0YukvRm98x/eBKVEcWUSYI5zq/kCIvzN9una9I41b85kI4sELv9DXG/XXGZQmB
WiD2TStBwVOGskbj5TE7cwbv/W53rDfNLK9HrmVgcmhbxGFihzs2hVjNbFeDHk7K
N0TWxNiPNQh2X8iJQ9sUAsI0a1XWoEaU1w6bIwjwUdCfVR5Qgw8Mz17QwdCI+baY
G6GKQ1r9pJFVwTnAu866CYCGFXcxkhwfOq0Rt0BWPy4AiogmQX1JxgPfUED2m2nz
LTJs7RSpcMTU30+WyPk6yM11kFsi0aEJ1TKslR26leLO13PmvB1DS8BHlPcfpHls
o5u270veo8erFkck6eOuk67iaoaW7IKJ0OecTEZKY/oJPqTdPlR1ODMZmaroaaeF
falMpWkUOuaPAfR51ajg73KCw697jlNU2/5SckBMbit0wgbQEIsVhzODKxyEiU6F
72H0V9XDmWSeyI2m8EUYGkSgnZ9glyXEqcX3euAByn9lDrZEydO/E0P+oPTufYJ+
gAs4WK/hCgyVV+aC9We/yk1upJUIQkoVqI0hDZVwhch1abZwxEt8/mJi6djp6rzn
nvdviMiOWNPelx8z7+L+ZRaLt2MwnW38qQwEhltgBiyfhwcC9gCGOpL0aRiMvbGK
WB2THQNXe3lUMptpYEgVAy+z4JIcGy1YONSxGEFLV7U3al4MmM2usL9eYhy2EwvU
FxN/4JMcA+XWcmkwWRH+QW7v3yyywZWbSwq5ddjDJ2JLqOOwIJPxAfjN0gGdg9bd
mH0SLJl8Bu2R8qsqb8XHNX5kwkZq+XDexwUk1J2RZBTzVftPZOiHvOsrjG8r/iks
VLWxHou9xd+s7CEohlv1hRB1IkCO53QXYVLGqPyWCDeiDGg9Li7hefSvH4baBkkh
U5XU18nc2Yt0CgeYi90HInPlXiBJVf69MwI2nX1CbDHv52MonUwBQDN+7tNgv9iL
hl5l7QxWgE9fn+Z3SVi/MdaNw0ryDK9JWN0kRoLLemnFgXzFPc2UdhUqRNyC6lo5
VkpHRXhJMcfzj6IBp/+g3c1u3Ck3NGSkcMPcr5EnYLvXkSNZq0xWWpd9xQ7bHpwM
iXyitY9pK6s7KtXCWLkhavIUGBm89n7ozMIFNCXMyhxz4rJDTQ0SjDn4/QyzAcr2
Mc0zP7FoA36kSAc5Y6w+Hnkmy0A3/ZZdBlcf76Nq/a+9JTFX+Xz00MESM7UIZajp
TFhfo2e4MHCCobHNHc/eqo5cKe4ijmaTy+aFAdc5Qny2HGGUDiwHjRj5zTRIGHTq
6rmk/cOXjXearr7KVLvwohavbcXz73cRuEtNOH1GKVnfjmJ3mrQPgJxgA4PXK9BA
C3T6sod6ypsPe6rNprVcTdRn7Y7c9Oz9BF6BilrSpKuGx6suZ3qU52suxBNMreQz
PVvM+ajdwFMj2G4959K1FXXdNvE9tDqGVRZBc3dX74t5CzETjyfC8O25z5lg5Si8
zJO4Ra/iK9+ufmLUW0375c7uIxEsf78Qwzyyxz19wqu7p/l8Vt7w7yovGHTxuI0d
4zlEHaETGg9vI5ogzcVR+RT3UQwi/+L6AFTIZYwfD0t6T70pRpcnwDQYCpt6h6dh
ia4gTt4ovHsmy3vNfAg63m9Ua8tm5iAdidCOcrIfZwMoKcnSW3ZW6yKdAyNKUeCT
I+loB6xtHsBP6rPtEERxo7II/CLcRILPtQA7q8HzaWAm/kmuwUryN4+qz2EyTWpG
uRyPe9YzqFjq/61nbkJg1nuyfhkrJTEltBqU0JDDF6kZfBJytrfIIFLmN0jVrmYq
2VA9j5L72VqVYh5k+ET6wcsRY0CXD05TrTieRQhGAT9DkKv5x9OZqJef/wyyEykZ
jIOrRrBKPdm1T0uy2dVugo3BCIB2RJwqgbNbl6gz5Ora1jjYMprYwk2Yb2P6+IJg
2RziGKfFta+rDV7h0u896pLlnh+ftNmryTSeEtsttRXsNVg/g4Vxe6beadBwbMoF
18ioFF7bgybO7uaYIhm4WYuiJ+vipjWhYVUBCP0NXmU54X+7LJt6FJAEVCX67nrj
FD7Yi0I1E+K7T/xfZ/HFCNoH1gjUzc2w32fhM6D4yohEFGAj/aMZXwpv0KW4h1VW
aH/LUE7pJBU2pU5yirA0nxe1N8dcLzh69Ec/o6gKyfNbBxvqOLBwU3ZWi/u93tyN
0WrJoY7nyJgJazMiS+q7bCFgGVxfVI6DaZ6twaP/cMluwI68Mzanb+XI9/Ay+7Mj
emuM9P/wew6WqBAhDTvgOEYlxcanYwaB+cWmhn7XKzHryUzkvP+fiCjaXtnLPH72
ogpB0Wtq6nQonXf6CRzDQuZpNRKODr/gULlY+iGzXsUH1QDPQrwBpvjvJKo0OOWk
is2nL/U939q7FaRAZRLVZowo1B+v59fdcmOym7/TqET+8ziy3kzKneFvFAwlbpDe
zyEPExgEf2MW3Dhbk5Iq5CjY0yoCmM6E6SsvLWivXQAwxGb0AwjA5POp+YPYs9cd
0KoT4H72Z4XaUQxQCmhqFAZPVHlHXNl2fUP8r/q1EUR3OS5dFMnDE1MOnPhOWvGz
TTEpFTn/7uvMuHvbqtDhbEJ9otQfwk7s1czNsOID9sEz/h/N7vaTcRXM3TQnhbJj
/01pIwmFDt2Iplbpj3JcPNF3qhTG4ShnQ0EEPmsKNp4CzgmBqJ91kkAEGMUTNCeZ
bAqhtIZA5oRXn7BE1+3bvzrNC5fEcFNujQjkBCnqAQr+0DzxIaHQfnoYcxJrKLTl
T/u/DCIznKCFRTThx2P1V/8Loe50DZPQ4ocOEpeMp3n3uwzMNHRm5FRN1CknyWR3
dA+ABpqmSeoPS56L9k/CO45PCvR5bLAV0UbrfRTm1aaFpA5V2ED+Xw2M+3Vk/LIs
9PpCojtuYLMWRxRz6Jdtw/GrJ3fHnx4kjy+Flq36mVKJD8ZWf/QaYyq3b2wii/y3
Pc3ySufNfYu94VAOWVH8NinYW+nq0IuXWHgwL0fZsfVJ05d9uGClQlL7+nLzMxhE
VZUN/lh0wMNUNuEvPxEze9MrpWaSv9jS6i/cYouuYgnceJ+8vO/01jV182RSCFBW
PLmRO97erbjUcXhH/slNSDNIiRUiACQsRJKHt++hLxlMT6CrgIZovRKFqmX5j/58
5AwPoo8mEjQ5u86oFQSaoK1ZjfCV9wrDQzj41wQiIAx53Ikxht6oGF86SrI0fefl
ZNiiP8WvRcSZCGgBWX1lRiysomWfLDROIw3/SkJ9c4cymrh4f50WQmftSLRZ57cg
nxsV0emydUPNI7DqTTQqEB0Vv+9sOaiUlPLXDYGCwMFy7+nXJ/7EDrCLKC0Zkssw
M+KaJ40cg3sBqPgzDUD1coO4x3DZUTVCtQ3Nq98vRDJyKI2cKel2s3dCeTkmFjkf
mGB1sP2aDni4YN2q1WSz3Jn61z+g9yMD/D5B/2GaMzud41db/YHcTvCVMXPdOy7h
nWoTgoc50WTylYjV8uy9cB/Igykvckag8jj734pKzlk1or3XyjTF+lcAQmx+6xg8
yL0yOuQ+3Oh+n7O9bINxdqEsjg463wbrNCDuaPCr1th5OtAQBjiTAAxjCszafuOF
n3+4tRAB/S4XAEofzsj5BNuCXJGRwVnHGS4ZOijpWUAJMhym732ccBJufLiMj8AR
aDJ1Ie2yzdF5+Yypm+5NyrybnnRYhcTupqr2qGcfhKfaLiMiizsjWI1itWhCCa4K
2FAekCso3IPYgnf2QpGO0qKEY2hE00ewpG8gw2Mp5yMgS5QVrwDMe7oVErMzvxoj
7hZieuLs6BJkkMvGQ2CbQQit2mhlP0kuF9lgzp3XY3JO7AQEH9EdHzs+LIWgaJFO
euZwuk1Nfh4zRZvsYW6PSouKD66pG3EcwWjvENtCUMT8JLnKM5uS6GUA6y3tlFl6
1wkgfaBSjrjgT0nyaRiqu7eDtSl/Osu5tCQ8aLrG9+eHn7nAK4pexLmM/h+5C9nL
oLuuPhviQkpqhyGO1LUIY4F9SNeMnOvfQlTLk4KSCiVejFiMdG2Lox2zej76lojT
1E8d1b14/GdY1DXO+61fqH3ca4QCqM9SydiVFA4O9nxEmUdRYMR+YYz9FCrPIqEG
s7JHljoNP7K6Bp2QKADLeTrV83SQ/7SeJFlr7S4VH/IYPiDa3UfXdNDDJs4V5Rgt
GzW7Th0/tO8ZLbJGSpQlYvap5zdBAu2nLM/ov/KcrF0QDOV+oOzPFNUhTaqxM+iE
XozqZ+SNFCspsPTSrKw30toUajOox4gXoLrGMr3f47ZSFC+VlVqGbdV2xDSF8+Hb
YuqHhaIXvPyRLnLDvHnDJOrD9C1fZJn4d5hVr0fwLt1fbP9paI38cCPb0kfvzJO2
R8oy5AkiFbLgtIpUUrHRiMGnpQ6ZSmfDqlIeHVRzniZI0b3f3OvO08nP/NLX0Gp+
hLUfQeTF9A8H6jVFiHfoY1Idiat1CpUFzZuYzmEyE958TlWrTb/gSecIn2jjFPwM
GcKM8+uqC5EAv+HGMyOTKo6W1dy97CbmEECuySJ57mLY6efJkHSGDAfAys/OCcsD
/Fzl3xYMzrGM01pJs7VtVD343Y0r9hqAcRLwG01cG646/wpysJmpyfq3Y/LXSDs/
eWeea5RaINTrdQFWXkxG1ZjNjPUIUKjbjL9JzI0v7SKPTprmeOsU4Bvm4I9HDvJV
Y2bgvyZlVuo4Ex1NORhZLPwPH80ea6Wo2fKpHajCQTtWfHhxr50NYqVxzASttbVr
3vWwXcGbZLi+Aq1Ed16IOgWEK7Jm2gDy6NlHgRy9wCNOBinzaaWielnfshYeWE0m
8US8qi71SSreL75aBT8eexuoyHbVRPNkumUm6ai1zfyuTdCCKNFirnpA8jYW5Ijs
lRMToN/AJdAPBvenoZwvRNbaAbAcUUMD8CLGvZ284Mwx/5QJsXXF7D1nlYppksQf
g3iFJU1bqwMn8nttwt/OKuf1KeZLdhfG+EyJGD0ZK3KtNmePLYNFSrDNffu0rivx
F5Me6Kzd79agX0BZPJWcLV4q9ALNMfog+PX/kF1p9Px0pIypRtNoTnpW1QVZALa9
/3f9Vf32hLIkoQrURpjNt9V5/mxcHyaKXcrTQyDit6mKhB2Nan8TE2Nr9AT1O02G
KSn2zcEjnqbeUBzkKNahdjMlLd4NdsFtY26fwCcmfK+Yw10XM4suhHv8Ju5ZMIKU
9eYxysuR1gV3w7DH8YQ+QJQHVDs/oLo61/Jdnysk1Iglo0KWAp4tFyVqf+CwsRym
BVq8d/duuq+Vqi01Gy38mhkayBQINqf+t5OgdebXQYAtNNREF0bbdsq9I2ha3hZg
9JlD8jTVIxpJxPGIKZnYoQttGCTGUI0ZiUvXhSlV04nTO7jAhy7wzFEIibvrEaWU
B9x3c+nzj6CS+GOO1ByQx8T4RZHctAHu8WxGTPNnOVz0A3F03Oo7JN/JX7wQQt3o
1D8VKU9AnqITvznvr8EbP1Jb1erXjMMs5WrnKsmwwtglJb671FSQO5d46+2OLOxJ
/Sd4kognIuIBn9u3348jZ30+TG1eX+0JCHsb16gvWrKBu7meDTKcECz/Zkos/7m+
PWzDZAQuaHTRHCL++ix8daSuePdAyFrmB5rmuDQbtGmThsanzcXu0O6zLT2gB/Q6
N8Nr2Tx4NLPMOf7XGjabVbyv3s1BjoSbTkQsmp9PF3tmaMc8ileHKRJtQqQY/A4x
jQ/VUihprFZ32EhJUP8zmzbg8f8+gCIRBEy3VajPIY5fyqzCtaOjTnZE/0B7iirW
tki6uSgHg5SjQ12D9f47ceWeY+1ckV2mjR46bVTdcC7kDjRapYgy5CTMmBFiyAVM
zgOJAbRsjIDZDeA01Ei9+d1qwDNFgcXcNyIGn9jzs+d8u3wYIlZhDcp5cufa0a8Y
UYCXSDzyJc9FNu+N+gbxX0J/tvagdHfzfg4yEXUMFAzuvxEbknvFhg70jtrD/zrx
Swn5fNvCxHOCr7BhVtXF9CNVdDZ/C5JbRYQq9shYVDAOojSh3xF+EzEEnbRZXaLP
RJLxDxFBNeAvXCabmv7tujYCSW0gy9+Nj5aXGCmkCe3Yiq1ZDMb+hLUVZweiCdyR
jN47WB7uIJ7RtiYXmw7BQzPwXRVR9H3+ZCqH+m1HszxO3TZIvBuApMMtL94J0zBq
U3idflMaMOjbUasnaxZaUyImGoLfeUSq2TznQJHQBwRUwij5xGqwEuXrOt2IbF5W
1RJvR5xuGpw3ALbYwNIlckC0BmQSYLd356EFCVyZyeazLHJm9Vvq/lPxbtFe4vah
6O+3xTR4DRw4+au5lQ6qXlDT/cs89MQen8AVLL2x1gFWY8H7TWHfFuE/GMWRJnOF
jnt+jHHtJ1Z8PS1+pfBajmwmsk71OCzOCl9tmyB1Lscd7x+IzUwUa7MORYNp8C9Z
DQYWyR8g1mGKN8tgM+kLujMS4w+xukIQNL+nonYwNKT/wVlGp7j/1Y3l1aeAE/0v
y2jURzApfNxMdLZFNkquTMetOuS2e20LbIc7caI9WC2U11tHOYssSbJRJSf4GH9d
K1OnFCi+DkQXLfVie3qHqCVA2WGaWFADuktHn67doGF5QpbW3x/KHiaLGANE69AD
5YDYgFX3KI5rYN/cXkVRHml1877Lgx8QiQ6DUU5BRBLU5nAcJ5X3Hyqxz/CpbaOs
yQVI9ZYruGxHY8fgdP/Ikn3D8VHnrGc6AI6IlINwEEV2wCyR4Xf7htkFx0Qpgslp
4LEQS0WhMVRw7Wi47GpSpLah3h5kl525lUxVLZkAklbdbFpqrK5iT7TIZUo8v5yG
wgggYs0KIqj+fGdXepMxMKFs77jshSRKb1tDnO8bezkU2KkfZQCj0JrbkKOdiNS5
gftL9TTFcgWLEQHttDb1z8zQorScmuJskgkh8t+Sh+q7v/36wCYLGMtvOjwHMdFN
I/1FHANdG8MVVhEW9ZGtCvSMoWwUt/aEOWVFa3n0b+Wg0OVuNkE0izcr+gZmVdhA
Si7pPXTAAn9Gk/UVEOTnF9oBY/5MT6PbbRvJHkG59SCzf5Cf8PkXQWd1u+EdA5aP
USzTE+1VV/9CtlkXMfXQVgEfFqCJJFHu10g4xORxQOvyURHCRcxBUnbI+TKG3MqT
465VixrolKdr8Gst8hJlDoEq8bBlT0oT6GVm5X8WvPEttkqVEI7Rk4Pylu3aNh3v
Le+PYjOhEqDI+9tD4n/8Las36nzRdDIiAFzxedD7DocrH3ufUuAQcyKW7D8V3Yyl
YxQ3n1b0Xgp7SUp22yncJzTm7kNCNUT/2DmVNp6A8JWa9k80p5z/vTgbZSf7S3AM
w76Znq8+wgVBGREnNlkQIW3eh/Zx+SqWFzRE2+ikd9bYC7pXvBu75idlc7eSPvhy
7QMitqQUqKSzbBa0j5tR/UUH4OOHM2VzncIug2dt3ooinxSvMMb1cegGTcgp7Cl6
EqOc0qGXd6V+Y33BNv7ECCWwAH0ne9/xOf8ByupfXOrMQZzHhWaHC6XdtjQK8hk2
0yFghDDht4DNH+jEMPnK8qd3wRXyjxIjT+/d2TnqLHfONyeVkL7w2Dul8CKy5/h5
Ibjo396Wxi6T8pSaAzOhfQRP/T8y1B8nZsHbPJ6u4OX0TcGsOUU5S+Roq2Llaqqd
r1inh7qOM29GU1h1E7pHPAuQPSZAjLV7yqr63lb+fHOk4QWn0mJ99driLugRn8mu
JDacJqujT6h1NDD9hlpabBj1G6tnwDLZ8CoX+8PdqgFzjIcGvAVQTJLJnnvk9OQ2
cdPuCfg7H+nwOo9kXXgwDYDAyuNOtJCyUOC0eQ+e11Uywb25gD+g5uxTPujHkG4h
vgNu5FFx88lvuVvtuRCwlNVAIgt5Zq+Pwtn571lswwS6lM3kFQMr+aFGE1b5duOf
LbXsk3baPTXMXB6MDytEl5gtRofrKLonJ9LWBWMAqKwrlceLDn4lMniZ+9TdaA5O
jhyy5954wNPm2fudyUuy8w6tUOa6hEXO9VbVrBvau5PnJGkPYMnLuX+Slt2zjIiu
OvqYK5/U20ZbQGqVf/E12HyZhuWeBzCsYgrtP9hfSVSvkdUQcKPRpfhi2XjWgPEC
S+u7zONXwOjWPq4o72W0bfK3OwL5G6rtx3ZkB9TNwrL6MSunFG/tXUKHyv+IJ0O1
ZFlZ9+7Y7n8XBlUJ0gIOT2jia8VsA0sK10/+nMBChalKyF3LENM8fbuH1uyVjjD9
bTzTHrSMjQ0HGp6OOqI6D/tqPZvyu2s3ycephpE4kgvTR7x8C76LdjYvxmGO8NKU
XbeQsrU9GYTVC3cj8BPGf0mpIYIWvNESNW5B0pnNT4dUr7jkHDLqanWzFhO+RfW/
sJpeSYSDUiVadYdRfzI54+vDCPqp/pShQH+8n0zZzI9WnSLtFZtsAp4BCyvim3Cd
hwV3a8PRQVa9wJGxyWOSLGU4gmnLYVA1HHAzXEvUs6KMNkSiGg5PLI+naN5MqX09
30+fWGcZNQEqIvueEmQ9t37Ri56wvBz4HK2nbhbtuzSth46JB+C6t++h5oQ0pMPb
I6TycrBIP91jiNZffKgCPT6U0vRPhmB4vZcu6NVgvcrbYwFqXT/nKzp5dLvtLkw5
aJhtgP6Hkm1Xbi8d8Krv8qXJmAKBJJF+lYYCPUelxxANHceGBy8RMjEGZEXRI6tO
5e3Q4m/oZ4gYU0TMCqzwmWv09mlyn0JV0N1cqMiGHqozuHn2BoN94fhCi6SFrwD+
e3Q3cFrJ/ZNd2Y8yTN1Qzbl0m3NfW8oHeZ2sJuRiASVNE0C/q7m4lem4m40c9rZP
KDGml0vuaLcUDI1pAeDiPeBFX+qaclcSnT8zxTTcShw1+CDUnhzspdufGjMhHqEj
+Ot2Ph07cuCx08bTm+WZoe+k3KbUVXYcJDDseLPaXm3q36snb7D5z1OVQX9eIu3/
JZEVt0E1Oi5QG8AnP8PaWm8+nDConE6/EIfZPz0ZAPFPVaLdT9Mt4HlrbBn0nxIX
7OjjkyZD+5fRZHK+x/JLUBMMwDaK0Gaw/DaKD9HU+WQ1RdgslF4YUu1Q+SL2a9MT
ORsazUPbUZiS3JEAr5021oKRQ+xyCmy0lzPenIipJonOM7x6xHDAepl4Mp8LotOp
+KfcGuRj8rwZE97VrPrfaBIa8ZgQ1UWjFUvRq5LO9tO6VUcyWXd0aXjqdugDmk+J
60KMQVmNqhorp6z/3WLe/xYm8OE9G4hYGTC5WGnDv9xeyqvOdWqPjpsRAE6jywrQ
zK3Q4gg2dfMdUN7WzWQb3rL6tDN7dJc1JMZO0L3zHNgcvDJQx90S5VBPEHq1TGwj
hCYw/Sr3aqaSLROkFVNwoKd3t/JIvTho9B4obK6XWNRduJd3pbyI8AQAKohoXYy0
jAao/z6F7o5JRfcUFRtAON+O1D+WBXC/3arpVRTka6zWpy4LYYvGpjOW1AEN/YEQ
/bjaIdjdlbH9gh51tL8bSD06Wj+zAtDCwkjCs0ZRfFEHJPcBE+kx/jzzk9oBRpGD
m10Hs5ioTCcH+xulQ1B8UqfMyOHwfEsiuw08IX8ndlUH4e6eDw3ICSuiseIaeLnC
Sgp0XB1cZe4gm5Tzy+vS/qk9/opOMD0BRJ0rrFDQB1BFP3E7++9j1zQQIPco1oQE
a7vijIv41HJlhAAHylZBhqMV4vAITbut/eag8feJw2DOiHrSpQWz3w3Zj9iyxU0+
Q6mEGI1xC7Tivs67fGpzJIMT1xjvEzSEDtZtZOdGSSW04DX/fDjfDoAcZLmYVt98
4PA6k2A5YoTQ2qgUTvDNrmftld344/2OE0OyYCLbkVFQBDXjwaehpukDOXKR02oP
DMV45nZlY4B9tZqExdL98tZuv21HHIqXlBoDt2rBWsL3A1iqeGjcBrjAjOQYWHgn
f8QWAWBt2yP71QtU+wnftcfXtxzyk+5hWGzVJynvShg3rv2TEY/KW6io0OUPsBEu
CqLxAQk56BO/8Pn9izmeqpowvXmhuwqBzXPLedBDXha0H1paqLB1Mxb57UNOsVA9
ib6TIFW1Zi8V2oksKrfZ3EbVUzlniEMyoC090QyyzGcnxeCkl2SULQqKgGB9oewf
M1Ubhvkf4/uvJmtcUvCYC/U6gPGyfIibZ2PPIxuAkYmNZdZ4sMNCIIJ4Y6DbEArY
+HWwpDHN/MEcTKHZqa8kUZRPREfTi8Dm+v6m81XbvRYGnYI2q706gwZjsfmEjYk8
ZTECpAgz3WZDAtQCdzEUHUJL4TM2HVy7lSDzVr3YCzyrAqJOM/kRMMnBQTcz/L9I
bFSK8H6OtpiY4/I7ZOOylzAWo4wsArqbJ2XkNqDqkRkf43jngMHuX9Z1m9eJkA5h
fH52TSGcqmCfhpUrkR5Z6WrrWAJAKuqvkCXTBXybNz0CCq+aX7q5NbsyX/g67aHU
jZYIUKk/Tmw2jFKGvN6ZIXRYerPyiVHoL/Hfz1PhbEtLhurWJ+7CRGOn1sJTwOUl
sdX2/lRpxOU09m1FgZRHJLLF1Z8MaXQhk9MlKhhKYiVXqvq1ZuVzpiKYtyt00s/C
Zsd2Vui84EqReQZNaMCIIodrvYzdjjzW6+NOe04bpbRvzotbeHr046M1Pe7y46bo
Cxt7naRlJRdlZWx/cUqaiOsAOmsuKxL7cyi9q/Y6I4VfZGuvTyb/jd5pcpwL6zFy
eldORiUKXTzm43geo29Nb67jD5HVM9v/01LDdbiqhiUBYd3kJjIsX78KaIHu1rG0
x3VAB3QcM599T9clxHTftKgJl0g7Xtj5kWd24g0R64RRjXn1D0mv7OsOax8mixRC
BL48xqz4j55mrl3DGppH0TkTZ7cQz0h4XzoL8/RR5gF9SMKOF7sBi6yg4zfe9kZ9
73N6L/K57Sh7070INOT+w5LdkdeppsWlYdZ6aOrIPIRYkkZ9lHZAFPSJrD44N2Hr
1vAhipGXQFlYtgnmwGtwMBVyeeuRKjGe6VVQyvMYXayqU7GT2NajQEraJN9qi7gE
zTzEEMGQeEaNlOKQEF1Mwj10sOTeFDZiq3ijYuMiAeRLxNvhr5hyeUtdPc4eoWVS
f4/1pvn99ybFuRoVlGSyGj8EluHukoTENhMpsorZObQ9RxrnfbeEgNWtlMQNdBOw
U4Ycw94TWnM3uBbwn0B2j254TqVKCfem1GsHJsOvZZyHpGB4uGD+Gc7QCEkV3OzI
xPPm5SuZ1Ch2FziNs6eFnP3a+oDJD89EjWFT3VboDyt+21Z1bnyd1xBu5n8vPK+N
xiwdcaNCk0Aley6cLufxct1HwWEMGyPjHmS7eaW/2sGSrB76JSvfXjqr43ejMjxQ
0rAzThtIOqD5ha4BzRZcM68eG3+WjQKhUX051W6cCsmw7XKLUcWv2eNOy1GN/Uj5
Agg9FzlO0uEGG9nF/IhMKSG4n/fisE1uxYPxtGo6p/VwEMj8BiOHtbLaneWxPvbk
tRCi1+/LR6JEjiFVbpCMFXtDu8oa7wMcjGFyLA2ks5JoxjXCH9j40Nhp1zgTPUnz
+PHXEWr7NbZJe29vdMUp6jsaa2gz+dp2qze8ZKE58I1q10EfIyoyuaXoeYe51jbC
QGiDRJYBC4IZlIkYy9q5ZaJrB5A0w0aEynlmzprWa3E52mHJrbf/h26vEST7eOmF
YSxfSh5atM+b87DYWV7gFe+Fg7o3OBn/okxACLu3+TRSeX2SLFyralQrr67PrAAa
DidRrv0HlLVZL3OLB3jKCGWw9xllW0xvoN6uEnklguN/FEyFyBmYsrxGlUAIdPX6
hotNJo+tXYAS0XMWt9cE8sECc0oywGOgf/NJ3fR3knxqD8Kg/y3MihwwomqOH8kv
X+OpUYiw6aUwHB6AyySUA0+SFazPisrLF104KxsMKMBWVzH6tznmYm6EHnHnFdz1
dpcC1GyTn1f7S4ZtnI18JTzcSi7Xh56ctEGbW56Gi6Evh9LH5YnoSSnjhlnfUi0x
xtuc43zIdpiK9IIpVK6wjOoss3Pi4JY6KlOQQoL69xre/6JTK22gM5Vce76xK6ZC
lGyPpfH18ulqAMswItYKCX55basnEh+GOx6r3rjRJ2AfKrR4/OR1QB8RVAcL/fim
6esBjnvEyXaUYZvsUn1Wdg+MFDcdfQy8F8patXWeD1pY2xTwvujbquthCnG2VQgh
Jeb9nzAO+TYJzFp/FmvMcbNt6GWioI8YJ5M5WWSzLjY6fcrfhRcQpHMopSZSZ9A1
JC982qmQBhzbH0ovOdiLQVXtPD2zcLx18GZCI7jUtq/mhskx2crtDBwJRiDRvEnN
ziuC5JHVLR9GTICs49Azy+SHsWEwn+s36lh5FMx5MM2No1FZ/TQk8qGJHjFu/hHw
2O2u2KLcXhzAFlQzD2miboulC9fnKZyCmqm15CaEWQqv4BhY4ZSJOpYb6sh1kJMs
6D+punePNjRX7lFRYVZcfW9WbmeMMYsaKQQ7ST+6yZ9TE3VoJp+7bhVlfIM6EXYS
8LgROuoXDV3saKZVnZ2xn9NKORQE+J8MtUtSWkWsqO50yNBCwvH5R7QJ8Q505FYY
Uww1oKqLby9bqFkFiPZteF7BTAVPKF8dCF2TU4aYlDMq1tErZVnbu2tOsYvh+NIQ
sWSNiOj4ETxmfW+eh5FcG6Tsxz9yLxCK7f+5Gg/c8x1BUHSf6eQ1E/28IFyV+1c9
RM3cn8oaG5/9H1Hg6/GUU6jeIfSQqhNeCx1k7d3au8VtLZgaxz8erOsk5hZ4oyNb
o4B7TQ+u1VQ+1rHa5ftldLlo/NbvN3m5xQ8FmfEMjdjTslsutJ89GNiiklyV478e
U9IBGbBH1HzG5hxWKG9kDTzr4hAoEdQ5kPYuHPRWjhbc30/cp49b/9fP4atASLj0
M4RJWq4Jd95GKnRLIPCYs14icSoC+dzNyNB5QjhuSBmdfk7ZElWCZfW7EfXGerZz
WT/Jj+u8qTVPjzcfeD6GtYPVZpxkPWkl+m5WXFH9PcgrjhU7AQ6I2KdopOf0T9XD
qmqU8oHl202yAG+u8rQI+loGx8sakd5UaRrqpTDPkysKDbjHuqCjFycG7e21fBgV
3+0/CTr2iAgkUQt4RHN15j/oeaK3ru8jh3WzpC4IEf5IfhEBElxR3SQDXuu73A5J
3ZWzZbVB6THfcniLEB/6i7w7hGAyl7i3xV2KFjTceQ8CQG+gldbov7H3urz6TRI1
A2BSZ4lwIk5iEpMuIxxHEso+zKD0oqNnWatW+mWkmrTngOPtrqsuz2mtaNiPVpr7
p0wBEFC8vQwxDo6S7xWHWP9OGorDhndyIOYL/KXG4ccBmW2rHuLMS8J0KzLSNrCp
O3vWgkMgaxh2TP5ZqNdIiX0qFMSxjddVP+13Ulmd8Z+zQay51jKWg9A35d5aVqPF
gv/r2LgV6GcvUR1Wqja/CrGq2HUceH5AKaOOA8hNEl37qv8y9jKgPzuiiDTjRgcy
ptuocYQWV3IcsWFi0YLrfK8pfHn/gbhLcyGNZzlzIlr/zZes5vWKVesC360Oma2N
BsZvM7ImVQpyXivupoUKWSJq/1Q76EHTb8/PeMfd9jVwZ60eyG7r7fSbTfSRfzL3
PV/ojO0i1YaLB7HqOx6BunWDd+jicSjO/e9yfpEEKCL506X8RuxuxvmmxR2FkHIe
QxzVpsG0XVgczR2whHXR5xn4GRhSOA7SaGvrabJOLBZnAZ+iJHZNtBicLkCfsqu3
/53wgETjpzgGxN7nsjFscJ6LaYix9MttETdk+U54n5X0V6s3GNQ3eiPfARQx5o82
Wq+YEkYULA6+fH9gMy2oN92Qpr6t11H0L8fSLoa5iD/wf0hovpr+WY4uk/8FBvXk
O7bthPd2pf9ozxyeyGaFs97gF6rOz2x8Odv5zog/KHWtKaVtj+BEQHPZfcm2pWLI
Iadfys+kBZELgsDx5lJWiuJrlHLVml3QdNtS9CYqqsp8bI5iPtuUX5vMj6EQZjup
qM6HaRQ5JTjBcqL5WlpD+ur17H2zWnC7IMCTsbW6lBBMMVaiV4EVzAzTG/Itx/BD
OMSwk32LQSRNrMcK4n5bI1E+PvL2Aca+qr/7dpYR4hq/1PdK4DfblGznqwOTgKax
I3j57Rzkpld/rx16S+m3oqhsCfIw0zuEAYIm1zVquRW0/KJ2kYheTE2E5Rkani/w
edqQa2OIxj5mvBPm8RC5rAMHAOcEpgnkTLXCB4vEmleY3aisYltyQ6vbIXZH6yAt
KJ1x9UiJECUl6bHAvUWOxzZmY+1hHW4BU4e3Vtr4iprq7USl5Ti7Ebv6rnxrk44I
q5HOwi1LUY15ay81h+nX7n/bgD5GKT5bsiVxgBpfAML+EFgcLCciGYHDBYosAVQT
3F0z5W16oNJophez3b0BC2ubAX9ptx7R1S3XKHn3V6jWX8bKIxApQkPtdbdjU4jp
T7OroH9Z4U9fIyblMzG/BgXc7iTMOodCfw4Dmo2/6PB7K7P1Zvfl0OrfBiT7jR3x
tvPOWz0+VPoCseHTQLwViqhO2M/9oD35CPMwplhXyIyS9ifdtszQd/30GNR8AGsj
E5BQ3K1IEXq/k9J4Qv5TWREEzqXy4FrvPGCwwoDm6KtLVhQpnBTdwX8ohf29W/QL
8T2ljalBB+lm3lvWsFGaPsRroJgODYxgHBMUp3DHrtZFaNl3d5R5GctmRgoq5g7x
A2daUj/JyGaD+tsGdn9FnwzeZywYfEPtDGiGzoXatffojM2pFI+3K+8u8z7JxGLE
e14Q2zxlq6gsiAecdMj0/yxvSRZHP1aoMXpXCEnPfGYfPgzmVsw//WieJsRltW7S
IfF+W36Aop1ZYRoX3lZsAdS+pJkYDmY29paw6hb1OAmbNbZLN/6qLpv+RcOXBfM+
aiRxaKhF1fC74GX/nI9SHvBoYomd3tAkVcxft5KA9hIW+0z33emgP9uDdFjJBk+2
TcTWdNatZve0hs6456Lw2Tnp+X0AWIi/QfC1izXvNyj4Iqv0BRlb3ArVKptC1Fy3
LEiJWjJHtSwW7LwHjsQTX9kyF4K42Pb10htN2329JPNl/HVu589Z2dw+cx4KilYG
Exkvk/OP09d3NVpDn0g5Nl83FkHt8YsZnQecGdSyaRXgepYEUJMTWaG02dHqv/Xw
dzbu810pXbDlthe1bbqYr51BkM1CRWP0XqItTuttM4UQofJeFyfdDgflXMYLyOS9
Ql2JxVo2i1WYH7BsVQsPjqT8ko2nYR5o9dHWLB3yJvxRSdd25Eqs/+SCSlzBX1CK
6ZWzu5evTlyU6JBNa4nwgzFiowq5yBOlo6OGzE16ZoqEE/nq0HbqSsE7752u5/9K
34yIUor27wwKCAegz6OnDH5uYEV0Kr9v82L+uxw6UlHKxTu1hhKs2wzKpVSY0l1K
SJuH72SL9WzUx953eNSw3WXrpn+pnaA0KQwu626qxPgKhVizI1bReuWG9XrTdxId
0KTDDVEbCu0DpRHrb+DbABxp7PiTLYisj5Y8mH0dB63ele6eQdrB0o3RLdk4C3/f
/j5gJEMpk6SvRMORcx1vK/FL9W9DtHNpxAW7mqNOfv8eUhhxHVx2fMogzaJpfsND
0M6nswFvqRkH0uaNl8ZB/V0dulie3shRfsE45xWSS7t+pVseJSSlYf65XUgSI2U5
eulKjNM5tx4LLcVjcKEcXXtZdp7UFQN7uZod6Zkkyoky0g73nwqeIIkAz8SUlp/t
my76PxYtop7xpAzmbVoQzkGJ+KXRlGYbzbimO1f8bFskX9uRuUbHV7mzlZ1+Rl29
odVtvjzSL4zJMFj2K7NQIAuy2HAMNg0qYxQUCuvdcujmEqoqujfHg/ejD0VbvH0o
vVsJlk5bSwpbZq77Fe8P+1CYBf9c2XHsOPxafK2rn7knAZ6p8lU68uYlqWVJDJSz
vCjCfoxQHRjaNtBaM8ahGjIKoZZ28H3+nrxKBpTTPDvztNJm5YPsWFJPF3yQvRGR
ZCxme/FAL5OB8L3INKFdqpNcE9K743senBplxM16zn3bdF7NOTMNNmOhyleZsQGe
9uW58gIsoelnCqT9CsuObxFGSPe82AkhNhnBxnTEQGYLvEj6PxPlu1Q3juIt/Sc3
r1ur81AwwI29Cp/luAbDYSI71a8sHcjR9Op1YwMCTQjHj2zjLYB/7KqVL+74TQUd
UH579blpteoIVJqwCGS+oJK182GRd+sVDRavRZ/5yWVRxwRr0FJVJ9EOG5c5zlFI
1BfZUEtagwqa13qmNOY/UgyB6anyRvM1vV9IJnSMbpdpZ46asXkEWQGTUJe3mP9w
OBCUU1w1Pzfx3PWKWw5L+5O4C6vCU+UfSs/lmuU2egDet17ZbQ/Brg0/nZGVXAgp
SmG5jQZpvQPVzAe8TZitSQ+iTJIxoGIpT+n5GegPUEyEMk5J7bSTYD4Umo8FOUtR
qGanXs9IwrOltjysJrOX2iRZg52tRV6AaRurVixNPZI0Uxa9Fh56PV9iCYOl6PUH
bwFmuH82w14XpFMt8pyFKumgjWuaIZ0b9JxRcQ9FeXybe2+q0QSrKUz5mMDmH1ME
j4t3M+hv3tVu9Un/DL40n99oT2tBV/9UTIDToDOl3D+kGd6l+cNYR7NVPGmrm4mI
rVNadGDsjXyRMSuFgMm+oCdrZSTxR6k/psMCRq1lvoFBKVAdptEbtxd+87VE0kYE
wAiJfxMcQh5CUBQES3PkENgnViGI10VbURpWcSL9ZO3sGlYFki4OU/zwgnnzuOqC
HKpR9704DpPTDDqmDU+7CxmrZNJ6EHdqEOt/dG+/+8dVFbuhaH44zLzvNR8RJHCm
ACOopKsf5Z7/IzXVrCc1EEGQCtaMnp4sFK2FtvZZvGyctmnOQdLwPutiyWxFR408
yVl1gwmK8eKgZsajOKIlx2Nuv2YB7ZkzTZdN1w0+0g26tZtTufKCFZ2ppyywFyq4
Rndp+DKLxxcMWTBEZYdFquAnJ43Nwc5YdNFucbQBRm9ZKu3t1TytOXRNzoX4lSHi
HLiKoj9ET1V3zHyYrl608EfwpApXpkn8CSjmrxFoqvp8401cRGhxtHlClTGXvES1
JKNOBahCUWmMcz7kqgwpXNvMI6Wbga3M9Jt8MgPOwznmraEvH2NgnJPDtbgf3+BC
G34xXhsmXd50dbichoduC/JTfn6CkHURu54k036edSQMdSuZDmxRx4mZyXkxsWIP
ZkZ0DvDjk9St0yt+oXSfari3te+JWmTTplg3fpf+K9fA1o6hbZiONBuM5kIx6pPl
/Alw11Of/voLa0FQE2/NzcrdqzwXNmj28kY7aUIM1ZK/lIfvxMO7zF4m8mNEGpHK
vAT/LlkST6IEgBi/Ypcc86fCxNhB1cxyOPY4z2Yh3/t4AQZfCqDK9rjtfD8qASay
s2jUB7kS3/Lh+igfELwqVNgVdalkvl6hfs6zQPK0eLHo4u/tr3oCvqBMDNkQCua1
p5Fzy+saxrOk7Cbzz6xov+GlWx3aqMkas2Xl25bPVY11twtIBvQG5IWIRdYOGThE
+1oZu/pPabNmlJmWnLtAE+Zhm8Qbnu6fX6AgD9pqr0hpYS1DVy2HZfJCfxTDF5+9
V67hXFAxCbzVphJyUFurbTk+VF9wbV1qtL/E69d8k/WHN85wfLqXw3mTgXZXSJC3
No8wutvfGNDhoYwnN1B3l0UaYfij+8uXOySxOngDr3H6BABhrOmjCdSN9NXeCXtN
ngWIAJA99tpFg9NGPTkqvSQD+yXMB6pmTbvSpMjm9BcyckDdrR9aT4XMHZzr+ytb
/I0bMSZH2zLXZTJlXyIZqpj+QBEXuHAFvDUPL4+VUjZHjLSnR8J34n2WoYvfyYau
s9lOCRGNwQt7vCoWqaBGYCLdYsH5qNnEi0XrYfSa/t2ax9sdXVkkBVPdj3SuXS79
GDwfQ67LfYayOk8fYkjDSTsDn5kF89WZTtJ7UGiMasi2mvUrhFYeOn6glZRiTvZw
09ZdprLMllcng4CQR1wBm9UiCW7Z9a/wUcUXSZyeZh/JFTvJyliw1Y3Za3xMnag+
U0Vo2BfOsGkLvdkA9qXwZF46uUAiBn0JsZPNZUnoIh2oXTVcMcmRmE0q7TYgoMwH
uiY6IMMQlVfvcZTDl4OGC1s7PtD9NTtlX3LOKKY8Rpv9NetfiDIaYtnPK5t6bt+L
MlQQga+TMSQm1i0WenNxNvT8zNEllxuUnvYQV1XdXEyrnCV7gHkiOqhKaFP/xVow
FArM7PDSUvfxvz79jRL/DKjd8Tvt61MPnc13BfQuq83eZtz4zv0kj2QdnFdYwsFR
2e9azEPtuCeqRsdd9U1ww5euOYy6euV5lNgshecWff66brQF5mN0u8AI2gX2JihK
iPWXNKjvSI/lVOO+w+qEpaXbqAq8dr7IozVzAxqgXQJdaaHdzDvRbGicHgeiSIHA
zV/M5dEy5CixQ11xp9XZP9/cOKmBkYPyeoNn2a9oCQC022Tpo0VqKhMKcLuaw0Wf
a5mu6qlm26zC/kMR49z64bumIDEeSipAi0C88eJiB6BVtkh0fU3CQVd/l+Kqwd+d
6shQN3QwOkrBnx6WlXY3KxAATvndIiZ9FK2zg+g0nXexVbXGd7KpAWeLjY+tuuYj
wa4ItujuUba+vLe6z0OMZxjc5Zf8qzV97O61vozvA9b+xkD6+rfhvzZLC5RHZTWZ
bOACJjBx+cV1FlQafWRJVqMKgX2NS06K9gKY4TRKXtB1cP3nw3F2kfcIDr5adqWi
1iBXo79POsKJnUqeMeT9uppk/yp44iC6dHppw52zYqyAWrjv82/5VWe5HSo/9kvU
9ECXdDpalhJSJDhRG95cfKIE2KZLiFGs9w3Taijf1Ug0DbRh7ZmOGcLUAf4POp8X
smE6cx1agYPtC0iS/q9K8fStSCB/XUJxXvCnwwNEalghNd6c8dLepQF+yZROrX0h
JCbi9tlg2V00vRUmPlf1Ls1RZsUNldsiHLcDAmZfG5isz56wO9L0cbEUX88vcPVS
PWXQIOn7pW9qrOWwCbJK6xlmrDsEAw7igbI0QJf1KlMF33kKXLVkR3Z1w520wEoJ
rxAQ8uzqHe2wD2sIlf7HyeU405blbayjEnxMEnqDQ73/wShyzJHIUsGNGvlyorj9
nA8pF1UJOq19+nqrSSa5tRVaAzBb5nvBtc+Ju+uwRryl2kIsQy5FBekktBRsHTcy
c8sP9eIeMqRAep37uMswuRUMz7j5V1BR1eijoc2tuRP1IxrbR5FShphB0NBKxYig
hB5QV3qqv+y1eNBLrx92c4aUVXMw0rGw8/xT/6PkylfbEYWfBVyg6mWqpIaffx66
uaKdCAjGf0EpFOYTtTGORfDes7hSa5Ijw9bGfsPa7a7gQKEBcQ/9P49XXyDI0q2v
U0L8OcaKvtw/up+ttdYDh+VEAWNRkOIaV3g3ZAp7m808ST86LlvY2xo2E61RHjbb
2Rh/5XKJuDonMVOKhoQ1Fz2RQh85uPS7u84H2RGKfp6VSibU4nskK5UWnfz8TJP4
SVonO719o4nQpYt5Ci9Fn1NpxcRNL9ilhvy4WPxSR2CxQpSpgymGhq6g9J4elX4A
dj46+DuIXEBURcwVfmAsgdDYKad38WaL3jDZR3jd4hukvsniUaMp942lrn0ATNNs
V0QIhKNeEAPnTvbcFlyfvul7zyYNaB6wHvBFAPlQ9lxTz/LTI3PjSc6XqqY9KAvb
Vf3OANGFanyIGx5Jp1PD6HtA5IWU9XF3GPxjMB+kUYqNvmAYzW2WR/pjoXl5q4YS
RA/biVjZMcLHs0eHFnGsEKSFu3+HLrGrV+0dKk23VVzGkDoK6IXSkF0gxnrSxqzC
gZbx7/Xt4FAPe7G/Q0ITCmpZmvTr+zIEVEXDU4PAPC1o6/DCDitlW1EYMr+6KKpy
/Q/aAGtG3Wz55+u1DA4olMNHvq4IdxSPkezdBTQQTbVsCUNW6216FWTYlJ17nhm8
5x4qy4fzvQo1jXqGKXeJ3l7pdVWPtmivhgQSkPHffLm/oPChXIIrnU5EhyaUHnv4
CjIkHc0Emil8IzXp/UjrtaEUtz2Ld+0rDLB/DK+b0fJ1+3YrduRcH/29/CWAfYhR
xYo++Eh48hmrOQxO1xtaXbAE+5HqDPUjWITSS82DEDQKlzmpXYQxLpkdwvOyihjN
IKPk7goRqchZXwKTAtPlwckfDkYC263uMylUFSVHFfNadOsC2hkT2V3mK3HButqF
UDGV1vyDsncQN5n4NpnG15fyGUfByr8flQCrDF4hdfEW+pJ3apDT0OlP4g0Dlnux
ZMwzhHGbkUBZFpZ4jcWmgSM0nDf4wr8AoI5U9W00sb/kXlAPxAVL2gSDNMXPuy6i
QvZmPFu1RKkNoLGrs5+35xALJocwb6s06AaQuvWdv8wS8Zf7zppYUF1Nof4IA9hL
GUbHzH/vORAJ/X8wFMbHQLDA1RGsm4C0L9SMI9R+UHqG5Y1Y4Pm3wWpAmf1dPG5j
d5J/tdUnQZQs+rMSXZIm/LK/r5u8lgEjKlYbGB5ResP+imORkh0+IH8Ru1ktdsDN
DirFANcRfaLbWzygsIadgF4RdwVny4JEV06DbI6F2zsLbe3MqhDH9tK0b74X1CmK
9vmcrxAwHDNkUWwNWuVFSmt+xeSUmerN/pQ0ZItFuEoh7b/N082fUcPuhOQTuV6R
ylc7bImjfjK5xg2lekxznWdt8mxFyYBARN5kyuNIWLiR07mhZFs4Hl2MNU25wIQv
sja9OI126+hZT0+j0Ot5WmYIWInNhe4mCUV5TRtByAojSfvW72hO4QZBioD9QY7w
dnmTNRf9lV+qmRDzUqZE+hl7rd4finZtxFw5MPBL58IaxBLy3TMqDEUsBGHXW9TT
ERq229pMPapn57z7+7Bx13FPMpa2EdCamVb7qz+TuMVfZVetHSW+NiZHIJQ14g3F
rSyPw6382IqJzYsMkUy70OZDIt6jTlTLrft8573/K5zNg7f+8myUtvyPw0FMLhkZ
1KmrVN/pTnVH27K//+eFrm8NO8P+L4yMFdjmNh9jYiObOAuo3dmgXErprwvsdunE
svExPUN1O8ORjtOAMT1Fra8o8cnpRIHZOMNMIRbHwO4wKx6vwznCBnVuw8P1Vh37
CcmG0BE+9bSKxFmoOY0N4lK2aXWfaYRm/l3RgS67qi+yKRXU56x1FxkpSJiemZMr
SV0lqIH3AXMASJV8qTYjtbEkr4T/p0OKVbsUyXQ2UyizU3n1zrHynPVkSXRuxcMp
REVi8D8K6SzzsBrmHgS/ZhRwo3CiBUoV4AZwS2JEazxhPiQFQUB/KtVuWfeXZvP1
S6xaZHOuZfq6q+1dV1frm+DO06sGaA+kiaop18hp+VL18ocJo0lKtl1SITC44RJg
OChDr+DGdP3ERTglxMWiO0UZ+Fp98EfhUy1edapAmFQdRZnq+I/oWKoM4vCxBTd+
LSosl028Tk9jD1YeeHRZpyrdZQ+eQ2k0ySu/n5btyxKZuKkGs+GCX3hbavk9l+Ga
XjlZeFM/fRdTzj32lF3XLhO4c6cYhuxDFCVYN9Xw7m90VvR/QEBvJiNnbRVnf59d
eKMBIEFOUCTVi7NwSUmauBrqTde8lDPR09oYMnsd4b4SPEP/GQbUSbkMddLIunVF
fAIDdSdq7FfRUJNaGmRLvSVxu9kd4KrqqLGrTdsubf2kRUSlFcr78ElT1+CSXVVE
MatPhK+wqXVE+jHAbmPgqVePE59DdHd4ZrM4gxoamzQQEeBntJxC+MuKKojkZLSa
uuRRtiBLRJ6XMCclf2pBa4W5sFtMNZ7HwOkNCQQy1oNZpwMJMiSP5rdzNY/kQoab
BtCyKB2+98WW2THd1NXEjVnStZ6C+hILqUYHWhDnC0M+WREOCaWnRVTBK8F4s2UU
78cJWDp8GrlxMTe4MKjJ4WV9jcONDLWb8N7tf1lyw9XCGdXM0fN2IeuvILIm5DXN
zUnPS6oms2D/XSmHLyIbrnSj1qSSG4UFYVBLhLcW2G5pGdazwLHaHFlQR7o0CjN6
a62tihh3wokyCZO0UY7Waq1w4sNaHIbc27jfdufkCeJEGVJB2/aXcfEw8bmpMCZb
5POfaIgihB12W5SeApymx62HapoD/0vi7+FdVFxIN541dXU4QtLpPVOGoA9eBJtH
SzaBFiXvI3dJT+4npR+qBofelFKmaEoAWhkYL1NLQMWxbojuD8X31xBi4Dagmuye
gyYg50veNk+vKNw45zWvJc2c4QKgpPeoC+XAyVPj0U/xpcRuBjbJ7SmFD122fj/J
FJiCkeaeG7P6eCF0XGeudJeuyQcL0UlXOtCIfw4lfC4og1Ihe+Ow73Hfcl71ugvV
6Ddx+AYk4gIj/uFOiN7mjzydPaESnWr4yKCwLYec9SAY5YC+dD3a2/NKfP0HKyP2
NBFSNqHGsw81sIb+HknJFbLLHjE0t0R0d0byCstHYrI3A5vMdL/oYv3dmwMJFQCA
6br9PJ7xTm67OtlkvuSzIjfHjOtEQVRNdUDXc91jVEZJey7kNyY4RuL9lMRTSdmO
EBSg75NIxcr1EWwYzdR/08W6L/xPvLdZEv8Ph4tHw/xMNpUHiATTRfTjicNwdDsN
VTElXdkNJaz+xyS918DwC7mQE7yTPX6ktT4gd+r78uA1qmuOhZxGLUCUqKDAfa3b
fqgPU4pabW+crKF6oZTkyfh5wzfFgFcU3U6PZJXSB8T3+92Bud813L9ChH75JlgC
C9FOLB+zhvutTFullJXZh/moihSLwocp1bbT+oqFePWpl9risYmjS8NF8zI05CuR
E7/jwavNZeHaid0UqS+7O1BJ80OMnTJwVM0yhUfEGhAXRiYMVuwsFhNRo+VjfR1z
irBd+TNTRDtPMqmPemRM9znTWnD+lfcaI/utIdl4mijTlOY71+yvzfA+smqCcQEw
4CxtubAbAoyia+OLaOlWUkb8TO7CqCcOr23v0PCX85TIjXVs52qk2EutMNAhnPxy
D0mnCo3tcl8ys+yJ9MSWXzUPrWGMcdhelqWaILrBBoxp8L++H+CauxSb0t+xCp2F
yQL6l9A/S7yxD7cdq3d+/dTX5qqFEMA6tLLziwuD9bW/aC+dM2nU/jwIKppW+dIt
fNnbFNVTWI8k07GiZWOnKl+2jyKrvsZMvMszfL2d6oeLtlQ8zJ87ptJyaSGjS4q1
Fz9/7SUNKxALffFyJ8joikNU/P7IPn1y6uTOvNGvYEmmzUGj+d43809Czy0mVXbw
4RVGcz5VPzXVUM8l15dGvUqIMGQbfF1vpIvNRPGsi3Jm/f/+MAn8HrgiasfRSpxJ
hVUQ4q/MqB894sneLTXefVm+XTFZLAAPyT8YgklauC8nsQSFgqS/fXXej2Wl8iR0
W3zygoVJlWqzeP7CWexrV6V9w4G6PB9tcI7VyxLEza9vOEzHHNmzRJw6iiHzEnO1
bjvlEBVXq1AVTi2XEBgJ/hSBMgy8J12+gAPbHtBs5O0eok35lakrw5RAnuJVB7c4
zLrqoeL6Q1CBs8UPULoJ12C0Hyk6SoAmzo6zC8A0P8ujwVG4XoByLtLzApv9E0P1
ctcPhgU4N2PN+veOR1UdrQEEl41Bwxqul2IEDaF4r03ZMnkacFOr/xv68/tfVZKa
Gzc/XTcHdBWKdslpJ8EH+0VDyKEBEy6MIXnZXFh3VMRay5HaBTZnv1Liw/0iyyWB
lKIZTzmvs/WKI7dy7952BDKgReexPx0Nlcr9MB2iUnJFUGuMYezvn7ZR+pWwHO7d
K31c4ZR0Lz4gSJOBz3oC8fnzETzQq0CHsVhBdshCgE5t/KYz3Wul2I8Ui65srVnp
6nOqaic/PxRH93ub+DRMDlll/6N6CKDsTnPD58jkQ7By/0IM0xn7envsVvuQhvL8
xkP66hcnHr4fFq2qho22JkT7ZAjjAOvTV3AJiYyrB0P8qzuDI7Ppw2Yfjo2bAbU0
P70weuYTpUOqyXNDfj/znUo7akb8wj4ZghjlUTHU+5Q811KuWCOdwFIPLY2NFB7d
UC9p1DsLV0HSU1xdxFZRPmzW2UGew5z+jlcUMS5CJEJaagWUZPkW5XiT8OOpO4uY
3Sg7DauGkTgELnfJIJteKtesAcclGj7AIHpziSUNWjj7FvmVbCwsG/Xw4C9mP2E2
AkIPF7mKEIMPDDgoiBStIbCqDKjXbxMz+ZXXwUvE9vEt4ldkfrFPV/XvcpsBo7HO
e4CYLBhoHqV8IxDlfqi3abcdqIf/AzBQ1AZFm0iDfqTD29QQMHe1OfhHKWL+At05
4km35gT0JouZJ5IGaArRn+U6GOGKkitghv6UT45SbFwMj0kYtMDTp4J2E6px15Jk
vD6w7x3YLAmQ+MaDmSG+YydJEPWWSyWlizGxe09ckbaFmsq1eJInk3+x14nBZX3w
4NEsg28bb9dfbSAEthzEOdeCkKjGCSfG46JRF4h6jqYu8gHvMIyst76XcpVwuqfe
xS6ODiKlLyqHSXXzN81o+NnySYVqumFbrmD9kEwJO1StB9GpuAP9N4jEw5BzgSt0
8LLfem9WaK/0nM9KcxJkn2V7MZuU+IyVJHYHtmh8eWiZPNP/zB5+kL8sEEULVwha
59Ez6t4HyRhp/lcMsCIS4ElXROAoZAaqdGrfpIoFItZSMHBIQIHgaVO4nHnYQUBu
MCBoyUtLt/vedvmW9DBMbUwsclKwnPtO8zrJ27bsfadZYlreIsKACLjre1SeDkCu
KNbrDqzNgORGGqX3R/IOEOT38lsg5BlaDhlfRf5ZOcsHpy5qx0mlXjumeeJeJUYU
jPm4st6gBp9zfl2FaelkW53m9Cdu/g+ecLHiiBy1+LAgSUSUNrww9FZpEB6rFlZs
ueuCGb8nY1ZAn6Ox8tacPDGUtl9T2pODymHgKsDEZMoGN1QYwgF9dBGoWbL/+kYQ
8yFbp8KJ1+2qJKxocwHvgah3BFZbT4ubjBbck10warBsKi3bfytDqx0hV6fbzuMA
bAFxZPfXvOuabsrNS4IfSkrHCIF/VzbJNDwrYUrteb/fL9YREurhb6tZLdE0GkVh
IMZe6f5rxk3sx0/En1AyRe+NVT3Sq7eBjqeA0TU+Jml8vQGest/S8gQKec3czSXE
/yOE2c51fKpXOjAszTSQeml828x97XA1HjeUPYeDi5HTgZV70452zvIz9yrOAQ47
0FyXOKE8pMalL9zKeF3gTGh4CnjucfoSGm8zALv+7FjdEq9s5uV0iGAt1quVgMaR
JHRdEAkHFln6NFvyJEvRb4x8uweN++9pk8CeHDud91+ov/D7ptMOsT1HweXDo/+r
cwmFQ8rX3t1/xpmeMZvNTpB5tnBLnwsuraJOQPU1cftRTvWPAHJH8ZEmv2JO0fHM
dJWwxFfPXVMwRcrTLE1AELa6t7xv+dgK3KjhFFcYfBNaNSTME56QxiOhLUn2GBXd
3Mtm+wLohBBhtjXC6/3flzrDwb/0dI7fooPscVtTC2ZHrI7RWpe2BOS2CqOLnj0H
EHbk6USvnY9wcLw3EMFGNFnEgwzKasJISEhYgFTytzFPP6r052FJxNph/WqwwyaP
yoAcaGk9x/sy+Nee6Ui7rnw+j2zcgHiEV+PGwXlHzLJ+DKQLuhDg9W48rYpJJqRb
pyD78JdI0dsB0oxjLGXL/hC/67U9dofv6DKDFcDUKVi4WlfEeTjll+ZFRILS+6i+
Ty0p8mV/bnN0mN5XJnbdrw5sIePVq/XSZZ9QII6M9FFSLIOBW/QOcVxF3UItpeFN
cnPCOR1I7NyEMv1xRskt9TuTd4vpLEyDTH3hDzCCH5SBcoZmaX9GMKGXqWlbTdEm
m3d5TTqjn2bOF8pZ0EuewQ8kOYXgVLOGVTBRVQACCqsl+4v5RM1xdj3U0mlcpcia
kkL6COqyjfd3393nlcb2jUIMfPdfoiqpB7xrOceRP0l++s1djsNXlSqaWgNfapoq
fu4RI0ruD0KQ7qrwk1WaeWswlnypPBF2l4XltHx/YQwjLRIQA1RHV595r4FRh4nV
Yb2MD5K2hEZsWaUhh6NTGjsY1Pjv6fvQ9KG/ZNGfg1jfUXqK72616fcYezZ1k3zp
xunCvJCodLIhv/jr6P61wOMwC+0LARqzVSbkliDszJBDytPpD2C70NR/XbrKfajd
9wlVEhjkHyJZ+EE0ymVzWh2OGAkAUEl/+seKKixkYwAmS0ZOKNAlR933q8Z9Cn5n
huCrbWr4vClmkHv/xeCWsoWdSAcsqJK8W5QJvsXAneTBXtu9R8F49O9ASr/0lsv3
Zp/jad/vWfdGmEPDxNqgQ0pH3HXhHehho5H0t0aejEhV8cEUBQtuKoikMk60RG/u
q794gVwLqJLX2CUrINzbklS9ojjDjVGePZb3akqz3peMP+41TROsw8NCw5ruzRCc
PpgxFRhDH3l7NPpQBE9vDR2k+5lSmcPChtzuGmvy23x+SImmBaLpZCGFL870IDD8
js0vqnCmqO4kZqHho76P09kiCwPU9JUsfVMTSbb1jCuVdNv+XxseNPn5vwu4xFqU
r0o2TiaD/L8kkkaB9UtNXWfZ5YMJSfIs3DCjhyXClv59hLdV28zw11T6dSnwKNyq
FnZsK3fSWnNd/6NxhQPQc8Z2/GRw4PYUoNUlxiz+FAIfFuIBQGF5xp58wrPE6PrC
NI3pr7zUNs+1FlgzyeKzV/y9G6RpWinsF+wouEOetUHT8CURwFr6990f6/OPdw2k
sKMvqBZheTUa2KJe9HRcXrvwGBDQAzBhfO8EOF5VSvV7QPNlALKrIKZ3/AnCezCc
jRrWVo9qxF6tsgjUnbVZ5GnVVTlcjoB/k2+RoiWo9DoGzlot7L6sTZMEDxa+J2HS
1lWU7ugfU6Pjo6cSdav7XJbOoJwy8qybI5ysvZBC5WWlRSFEU6m7sebXbFUrlCyI
Q9ckQFI0/Z5nZXsigY+UHH87GE9b/OdP2Fm0c/jOJXsRqUSvV7RqlxP4tkudxgcX
SK6PyST0CxkG0yLDZqlLfBjNxs21a2kM0QCMfZopuaPZ4lE94TD/xoehi+o5PqHf
fuTcCgxV7NVaKKEWRSIGeq8IL3DToEHjTjodTx3/PXnbi0BTDa0ZYSS/fxdca5RK
HX2aeECouoaCw0hoWBFPWX8UbNlpMmMonLx8phC8UZba6qiugxrtb3YqdG+wo03U
UEGX+unmJJ1AWN1hqk4shj6zj+gYCDGaTp9nQyLEgqW8+CWleFCgMMe6eEuEVBq+
WxhG+CQzqbTv8d65c928563fElYlkMtru7Asn/jnyW0xSlwnrgxsE+CGzrh8ND8n
Z3rrB5r/76V24+S48cVWajb/pmlmlsFYD9mQE+NNQAhEIrQNUFj5OeUOUHPB4tSI
kXZBqmri0dT3sZuD3sEw1b4cpbSSUyUpVbSJlktRryY4CqN4AmJL621CTPTFClF9
PtXEZMHvBseTc7KNVub63MCCx3qHHEFxxpjGg6DzLrofbQT3WO1Dif/7R/CXfDKd
Wr8QlOgk6u+V5pA2vLUcPIItzsJapSK/ECbYrAyNxc/3eWKn0Edb8ViIXMigZi+E
m4f8ea2kFvrvNRzMdy9LHVpARnf6UV+QZOWeWe4UErbNl9/khfC2xcQatgRPjHp5
QmhmvAAT+EldaHf1uqDjkc6cmKBUZ3kn508SpGAR0mMW1Fub1WvqZFZ9MnaF2Ym0
6yrvtXsWWf4IxmCQkNwpNRBMdknXFgbKGOtJKTl39OFfibYJ538d7I6K6qVDZC8C
aXDIjoEKm9J6AwV3BUubzRNIWHphplWr6cQodOsHzmssQKSsHPkcW8/xIve+trEw
xEQeka7xA4EgUjQj/KcBo+/7FRvWIYC0cX5bbL4GUYpKVuUK+Ak3xcuH/BUhXEdC
LJrQ1wLPHyZEo7ZkTGtJIdEvCe4yRqtqz3bBFZSPhlL7X9W1Yfoe+aMi9akwavZ0
CsmfPueL3gnDvnKQlse+OAwL02T/byJYTan3AvUXa5tJ81/cvBNsp+MH585Iwcpp
XrN6P7BVBd5wI4/uw+iVYuxLoEbcOM1Fv+50xSZLrIGmL7Mlqg2X/R1tmmSliXJW
kT80DInU1VQBDo2WQ4t0LBI1AT0399d47CS6p+JR4wAX54Y7GJO5lbDryNLmq4J2
KSrxcfqKndM+ETRwZAFtd/EC0rzbxkxyZ6BdQTJxyaasTi2hE14PstpMYPJG47RN
V6RrHBymOeB940hs+VTVlG+4MX1sGEo8P0slJeLjffCRoqBwF8duiosE/Pm6eO25
IvtuqNgrW/ypSD8E5173KbrUzB8/SNk5tE3wCP7KW9dRbFy6s23LRXel1MJmJ9NT
22gxaTy8g0xguo3zO2GpME4cWU1wygMjBYIU1Bx+QrA2mKwJ3bxJ197+w+zGoP8a
JU88ZcDollvmJAnSnfsaUV+3W5Xl1TB6d49vRcUFQWyM+bcJ01E+4tVTjIuAhQ+f
VwNkObI/uE2DAgL8jMWoVRt587Lx7sxjSYxepxC5o0k/U3j+AeNA/76oMSjwhov6
Yuha0ewkGK+9HLHb76IuHKe+dtfOYkKGMHE4Ji2skZa+HxHf+looxMNqaIjJJxXj
WBldX897uM0ARy8iiABILjjkERIB4PN6f+VALGD44kS7X2yU91tVVgxpMMY/2lU/
A71jO2luneiRc0bEBn6TeW+sC/BMCifZEGMdo5UtWSS8oMP5TLR1UZZt0MU9h1R8
aJj7yRPU7NFZvf4cEUN/HiEgWwoHWBGDYDlnBoSZi8f/tJg0yTZAKO17lHDrQIQX
V+7Zye5VK+oxTjUpX1G8D66DJ9rjE9Z5M3GFWu03V3UegxLd+voYyQq+0/MRI4UU
KAxP8EVvbIRYLCcdh+0kK5YhVkyHeojqNi04oqTmmqLmjJPlEmm0oOaUHCdNfmx3
60UUrZKrmlRs4ByPnKjYPb5wCCTadXbKzqLYxZW9fQTDN3AQIWBPYMV8WzfYYJfN
Cx8lmQLwU8EnLFJ6Gd/KVcPfO1z5Gs5jZ7m75LjwI9qrSYGyar/gTDknvYkSNRwv
rap+rhddf5DEuuo/+TTrCk9CYnLq3L4yQmkM/a5/+5qeHO2fI8qg9X2+fOKLebPd
M8eMnpNO4zxLiqkEI4EWSDDbaeTAe/xG9EgR8QULO9I6iqnZPh7xX9c1lVFgXHCj
5lfKOpkbMozhYBcuWypgL5YvjKO6ZAPLv/ixIk2GTFPUlGpZjOrL1EBjkAs+rSIl
KD+Q9wQqSIHcHuVYqtZXxOs/1ktg93Ye/HZBkmuH8/875+cOPcfBL58Rp05Zg0eM
YrOJPSFgpLjilY/S0V+QqxloN5okKvrJzZYycJWKN4BCK+kZBOnifZTsD9iJjxHn
sX6Dka+LnLpu6HvjA1orwFM9mekUMsqAnbxjHpiDkvjitxCgGBPXEdnCD0wMu9Fb
vEtU5MYu6JBj53NHMGj0XhPgckSP4Y71KNXEFbnUnKKUUOZapIUDQ0F3YaCOwlOU
dMsLZ6ugeBPw7qTdbpNF0VeiLB/zXA6tB9a3PW8ABEMAvUFxtmUuMHtCbvDl/j/Q
noVMlv5qSUB2at5L3EmXM+RrbkfmiuBS4txYxYmCqYQmFUWjPXBpyJRQXn/HLKW3
ssJ2JsBXBmOEJO+kJJSo1t43i6XotMt1PZPtoatNLlVMLeSUgD+auXZFbbL/5YWM
lCv+oclP/d5XxPTsGY+gc12Dkdgjc0MQ352xBKH/5pqYLUFEsE9EMYSi0upxpUNl
zMoihm3zbrK8rGizTaY3IVeYeRxIsPxQIfXdukv6sMoWLvew/OThYf0GWoSfB8lQ
lRBcyHtYru+lnVB4qv1EFoG/Iu1wU/B1WfCCJmFZ0goUBQ0oUD4X+jobwe04L7U2
XKKEdkEnbuTkSkmFkARaAcbzZEoPuLvIDD8wp9gToxbLitKFL0yoBKz0ghZzWvoA
Ta+etXCcFEDUHDx/Rs8Mf8xEfF7dgvfHGvO6Inai73gnz0+atB9CeYObKMTEKYE2
6t57tUajRC0l7iBH7uCfXQWfc93QTtMBlEAeSZSvymvR+X+4pIroWtf3ryZlcGCX
eBPpf+MA74WeI9jeC7cJsvB9TwL3U6QmbsWA6l7h9Re3yF08QmqkfOsdjAQ0qT4I
/UXzRVlprRPJEPO5VbS2lnd6rObPSBGcmxUWW07ULWGhyPuhjRA/ietM0vFWbi0y
zffUMOJvf0cIhF+9gJy5L2uAyUs6Eid6Coof+1gw9ofnjQhvhadGA+9dLc64SFLf
BqpefApvGkgHB8kA8CsT78WOgPZhwjXzB10LJD1e0L6Y423h7XTYngFictwF1743
gPVR/NtBEptrYtj1NhtgohGGVLhtGNV1WyfUBLK16QL3aWOCZ7lOX1WrlNUnNU9W
ULPZPNgR9emf3LeoLfc+L+u9dAa7T1bC5qRHkipw6uYvCEFA4Sdf5ZuHAPZmlCQH
bbyfJXjnqd0Pkk2lJLGGcKwv9zdipW2ztMvG9KybTeSXW8dlKNUimPQNNe/L5IuL
RkA0kOPs3vbF8Zk5QS57L6jhMzIhvpRkWRFPWr4ww6ggFmhsVslCr6EeNunx9zQ0
/mUS9/4mz4ZvaxBXhrNRj8XCrJJTyPITfEbe88w6oA5QuFHHR5WKosy8aOFxzr1e
ImGY8FPBnmcYHasGjZfNDjQJYbyp1MXKTSgDLfdsEkgsC414GRSo57vgFYiYdrE+
iJ+MvZLoj4mNzAn85KYntay/qJYDG3v74Ogoq4XlH0JlBEgB7f5DHB1Ud3QiZP65
C4G+UVCTGXy/2908WqtFs955A597ryPYyl0s34eCEEXJXQqaohpSb8U/41MxFkpM
If7BWnk2GM81t9f1YtxPIlQ+AAaTaTQ6V0AYyMnWQqlEm5UF3IwIMYWe00/g+zil
Lmdy6f1+ZMKUG7ESwHr+Vg/H29mawzuSNK413DXd1MVulEWh6VrEjcZSiS+m9mZB
rRMtBUX6r4BUrdatEiJNwLbsSX3EKxR1sd9CtFn87xl+lkZ0I2+5LgpVwHztld5I
yNGOnM1S/YludNwWJonNKDpLbIHMeJrEcqzc0QHRdkKQ4ewxD1/sBsTayquK3MXm
/kgelMZ4sDZdgcDrAtT3aXMWspHRAedl2NMlfiizHxqZCqeFekqrw91rtNGZgvFy
bdsqQ4M+2zj4wpuTAguwCgWjn+YyNcrhy0pIz/pd92AynSezs26u110ZnjHaPfzF
t2AjStzaAThK3dobul5B1rYfujWT1iFSofF/dxAC/0tJc/1svF9N9YG0oEuFJpUG
oDOra9UhU96HiS6nP0YKdZnOK5ByR4l2qXwGaySlqHjttCbKVsIZ5GY2JICkCoDf
fRWomhaR99xsjdHDHBXfXoFdQ0DQMcc/hJIXnqoEfdE/jGD79OR/usMY/vAQyZT/
Um1rcul+j0FoTwtFbT5U3upe56VHTcY721n4V4C72w1Lr0lfwZCtvbubcWAyHGX6
GAdXIKzU1wT4jy2Qd7t68kb8MSZPi6RzBgvyy91OOgeBjyYXEY/hor/MWwB58iEw
sRwz1TKgMbwFvcOD8N/uqrnfnZtqy3DXm/xKgDrcOEz0adlx4Ih8GyVyJykCRHhb
hTgt3FBCSV7ZwCPV63Z/8H9amywk4dB5tgOdR+f3rXW/wbPTorEShhhhQrET41QA
GLtNfXqHYf6uY0UdvjmSv7Y7d9lU1WPWJuA97TZ2/Nx1NEmEyWzw9+nehoKbtCej
KdQec197Rm/Ki674UpfNx2ZsP+j3uhMAOOSephYUMr/zCYpAqxEnso4lqyY/sRRU
yUZpiFtJGqbsy3xQkGvJ/YHIAJQvCwuRT4XldjezTKkCXDtvNF2HLH/4Cq8MxVf/
YH/PR5ug07IuD6G5WutC4UXFj9mkbbBP1n1bqOya+XJcG1HamHihN2sA1trhOYes
0ktIzWftN9AiiGsdPcmopYRdWsX7RdP0KIUbQOHHGkReLmpmzAS3ZopfwwSBvXPg
zV0bMXA9TjWx0yrcxLZ7ihSDlMlP/yGXvETUBUWzKAZ81VF1LRso6I4U2eNP6K9E
BzqKmOnsbtoNkmmb6HMgZ7ZMaa5WkTgsra7ePik3Uhf47qEGz4vRVKLd7TnMcrz1
6rcQplj5+nGqvvTAMv6UEwHZceebUXWe++B8qLSVvFnofnjqpL4Tsrr2R0ADv50f
StyFsb5K606s73tH3q1lC46B+YDmo/J55fnyDrzFetWFPaqzC0m4JT9W4/GBap7U
k4BzCTzccSc6CoEWVIFHyw/GdNW2ABwPGY+L95xPATZkx6HgoC6tkX+2xsuTdip8
UY44FNHbPVKsP5/37oZRtvpPWuyS9gz+m5p1zCKgCBSieLk66TavQcHdVEbgJ+NJ
HruVfXZVlV1OlrCNdU2hN+GI0/MKB7SrW9ic/toAUN6xvpLddPCcE0NVYX0JpQTU
R88Cu+5rfES/3rZOZtLCaB5wlGTENMBZxEKKk/syeelrUX2Ukltul6fnbxSjlJNh
xRYY2h8Vq14CNer4KmJLhdF0NjKQ9e/mC7uikYiyiCNfU5sSNAyLl8PVEo3cMzv7
6tb0LpbFr4BqMvfiLi20NL0MqB1x5R7KGIlw6LP9XKgpktyzelKbMeDEr3E9p98a
URmyoVBzIkoioFVZBv+D2tawmH3ljZU/GsSKKBqwW6kSTNL5l1t3cCR2lqTYKg2f
dE75CgUOQAsuuADQf2id6vglDoCw1gN4xOLFloS5G2t+DE7N8EKG2z5iafkPMz6o
1FyFQNkWNTKKFyyWkymXtMZVPyR0+xtwRWaaaBA8q1OBApRfEQUHTDwdCiSpBxiX
rahsbSTzJg61qgl8v8GPOKOYXwTvavvLFfI8F6ugXwMl45llRY3sz19H8Lqpnwac
CBsvy2KRs7RSQPk0yfPSg+zXvO5j9ykZcsPwyBmfXLVt7pQTFHDixZRtDtiXAfl8
VJU1HLZKrPkrz7yiuZCceLJjRX5vhLEJaG8D9ZvQXSJyZENTxwxH58Xm6n9uXKli
AlGaoaN0xg5IGJI4pmngBmSU1vCoVtPUj7Gt4odFR7GAWNb5UtqjDNgLXq8bB0H6
mCIXhYW8Q2IcJlXrZiONNjik1AWQxiPrFMdhV5nXae1mSSxBgvMQUsJEDH6z+ZTs
vCZhX/+yY0ILPUE+/CKs+jgP6TBmP58BQFMsMqZULLja6TktVkwnrtEg2ZvX8JLS
oQxn01vftRef1RBD4eHW5lhbclzSfBXagOagPFd6A8QLxUqRrcgbM3+zAmYDO21g
AQQ+89oCJE856vAGch3ZMyaY/sV1o9OdzAqsMNOg6nGcpIKcp+9Zz4tNekFNs7hE
9yJtCfa/PgcDPZoDdsfm+rmLZYyKcAfom5yBE/V947sKjuW/qxGObIr3ax+rYK7Q
sUadO5Ep5nRVMRhafdoGXSyYN0QuWK2HtykK56OQpItMRvFJta8TNRO5bK0MCEuq
w3t8YBErqRdwZ/MnMrgRjYWsYxEqzrHFXAGWK+UvbfONA97uRNC5NAu5SoknKTtW
Gj8yov1MJrso2vZYvFG5HN47ZGhRaWTSo5Zh3xENPnflEaj0BTupDGAjYhAxhEM+
EBG7ougwJCOgZh2KLjW4moSREMBSCkXvDXh1mow6J4I0ufYilSCib4snxiQm6tqC
oxHxOQY2T0HhoASMwGMTjXjhqrI1WTefhYZoWppMtaJxaO8+q70+yTtEaf/43tdB
AAn9ziCaSGWS6GM7+flTJ6h/+rkHd+mi2ccp3NOeE/OBGSnmsf9ZBTtVrUjhVkWS
s8VsaEE1QxoJoaXYAFchZh1g6Dc2vJBVIPpIBm7EFfmHWlc1l4VWMXfiYInB0/Ln
rNXYhkgO44v2G0ofVJBbZfGuEnIUN+dapNqTol37a3EGkxgJfccx5e5FkvNM9da6
aOz0sMr+MsdznKf101Xh9eci6oPZuSC6YvZ3sE0I7AmH9iF6v0ZKSyfcxpJ1Fhol
kjdMwsavNWrkaTVhH4or3DwNQjyezkVkVhkOm7qybImULLJOlBmfvi3gevi9k/7q
brr7aWHYGpJtNl2SM9G2IyoZEYVdjeUYEMEMXna27+iFZtMtsHZpk0QUsxsYRf8O
sxUs4CYQ4asTX6ydPR3GLCy5b1TTkeGU2O+q15ruBH0JyTqqPKGejFoUlJB0MMmr
8Di+vxgH4GPfbkRderWJnnK+ytIDT64+RtbgBvuJ1+bxPcqhOZjtSnMhvuthA5Cm
OBwsCc8ab39jrNJ76ydYcqKtLXO98kpfV/ze6aioW06O0j4j6zk7O3rTZFxWcN0T
sRK0D2X7kjB84Oow9a32SkLp3lDBSpjJ7TooVokysuH9n12Ho4dROVK5uGm0mH50
FsdTSJcrS3j3xWgOXc381lLdM9HMiADFmb81OwKYk6ugOAHPRBBhmEyQfg9fPFgt
B+A4i7eC9V4aJuNDnCS4zoVJya/njZH2cXHepaWg2xedN2v1G/h0ByE+Qa9PLe0a
fEV6VndvL7cU1yfYfGjwcBuHOcSjC7JfglauNCKFhSJK0tDFI32PE327JHb2kyK4
TYX7/8/sdtw2WOWMyPslRFP6v4Ee0SZi2ha+Qj3B2K8Kp1Zizt/N6CNjWObBA3sI
kzXEATRE8tAzAJINBSUtBXthxF3evCH9RVlv/oj2+tXhdcmS2GbfwkExs8hjByN+
y7khikMp3EX+uAkNsqtWWOgQUOEHFrjlRz7yeOG/eqjtFL37zwVV6llM19a3zs1D
gedO94KvABLNS7/cc+ABy34/ZlgrzzY0zNPuxlW0fudUCwQGWKo0NUE8lwVcH/7W
C5yXIKDbKpbBdnAaTGy62UYUDvXzhcMyaLdJGLjU/FtNTbo2V611d8FuBRrg9f7f
X93BmDe1d7YaDJ9Ytb5FpeKRLakAUYy07wgQttFqyWC7mVUNPls0oCUHcyb2xUhL
AkpM20XSRR4wgHP4Vrm4VKNkOcOy/t6E85RGNtQWSKrt0qPToBgCCvgHu2CYadez
s31ovbc3ztydXxUHbQ/vYjFwzkg5vKKO7pc/ezV3rwG7ZIlI3mxpFugbubWYbQ7g
yWBvSsgwpYsfUxvcc5WPQknBq+Lhu7WHJo4zOYSbcXvVb5vh2xgFFAhEkTOMN8kD
XjDcbEFugnYjkP0A03BcqG4yxwWPIK0v8fW53J2ld3H45vYTIASxPfMauhPTSnGv
66mlCWp9AniCcZ6/VQAXxYzvxFLuWB4IGB1c9G+2n/sfpU1OIGORRrKYFjwNDuh9
KTYxVsnTcTLsFOkPNRiIsH8xSuaowoSveWgOWgcMX89ufiXLYNtYkmxDsrQ+FfKa
o0hWbG2kXlbdCot0uybttJGFAfn5x8JqgSI5v7D74smNiLLvhRZKWcwnuyBD2XBu
pimQkUpOS5u1huOVybNnbf5J42g+9k+BgWo00cCl9pLSBJ1TqdBO0526FA58N1p2
7lndBDaqZDJqJqCf8wUHfqPyV0Imrc4CwAPgYmty3N8wVpQQfMpxb6qJxjRVKl1d
iom5i3ivXheUkDkmAZOXE+Z2SdDAI1Le/vNgCo6EEzfRvIMphjXj0sdpt8ZgTsu/
zIQhw++WoetWNgdaPp6gJIE9JtaA1lXhTS9Ayjfw/uRA+Nlrpsh4UDUy4YrD6tat
Y2biJ6376t8Pf8f/V5VQErST0pcyp6/UcbruqxUIYfvWnKq5grsLTZurZ7xGYhqI
0R1bKBdvadnzHASgBWJaxGBTvSW8mW5OO78GHGW569JwvRRIiH645fFA/HbulBwu
sMZdxPXNJLNV2gwRlyQfnxNg1BcECcpFky+wspwhpNGx4KmnJZpzyIGOmN1MqxTB
EZIZAw55PYH3Yyogv7Wdt6KaU3OHFClpVL5rMIZPyg7uSLpUo9QtWzA5luEkonLv
tOY1CjuFhdgHCaWQxLLwFXvluFoCTX75wtUvvuAgmDs3aHCC9WgD1qlTwanNwuDr
yvQ+DlL6ZiZ4hnW3tizYUOeFJQXexC9FnOS9rFWBJLmvmCWluqnTFAXkCfi51yDK
8FND7nH7JwFV91KtDD0l6BbtIYQmW6rRxCW2T+krOWjUTSFaecy++lStUQnCdCHM
Y3Weg9LLKNhTaqefF+3Cz68U4323Fg1CM0WBkp4nCBMi+/v2YTpRgsYhzZp35Soq
KaM5gQe0RsNUp94Yo12+HfJ1Gbp6JP5s8cXAkW6Beapf00FRcVejSRrpLTxNr5tV
R7QZ+iBFds8GAi32PvDNzeVXAAFsG1Z8yeo8AuBWRLRyRVLCcgnjKdgRz1NaIWkI
jN34lhwVNeBbjuMuK7C5M/ejUWvzB7bTnJSqJ7lQfrPdjzhJyA8qH40uKwNwmx24
mITY4MQOrXmyzcEx6+XQZrBtb3k0+hyMzlZ8lSjxK/sYhqCF/5fETCm4jUiD9a81
LTBTI5pAcUUqS/ikzuGONza7DpNRPF51wMzQGh5icOjcAtOHHAPFgO0OVHgROuCd
TzzeLVsNhcOIL5MeF4GvlWdgY5bQyE0aEzPzpR9JQoJCh9bkxRcKAwxUdU35G1Vo
Y2/KPDjQ0UFsSLLrqh057GWkJn4eQT+iLGkLg+xVSSBPaLQwbDyu/qOyYDrC64PE
55jw9kCVRWPHqmQd6s32ErgT650uMaT5sv5Ex6IGsGQbt2a8OSHzDnhvg/DtlfH1
6ALuwcrTYc8x/gGft8AlDEoSy9RQ3yl8cHH4BcASu3pfVDhNR08OH6NqvkL0x10r
U7hylFymfEmRlQuQsZuxam3z+nXfVVnvhay4brp9i/1XdWO+oA3i7ItimDXVNi39
vbRRHzN5B0gCKn0dnK+3XCI3RkxJJJUKTc2UcFbczDXJS/YuXBgSWtV3OmLIOCzJ
vS3qDvZuxtEPJtJ0FXqBnHvW4pVgui149RHZtSrKPbOOgmreecPMzV1H1v2LCRtd
V/r37Rq1vWY5Dd49PhuwM/y1B5DRfqKbeG+zF5sXB9jHRrVydwHCyOyVIoFFFXQg
0zG3VRjAHLAICRUewtCD19hCQ1juflf3N/my91kpIRJNxW5iqtOcaFqowq0s9Zgz
bLJhugnrZ9H9q93luwPwzxaycviKSk1vyz30WWpKpARWcg0USN7hWJ1M2gKPKz/1
CD8PI5QcffsVCsUwrJRx4dfIPtUhvqpw5tWCKLWkzO2J0qTQBGzjxUhrigKohyWM
o9A1CttXlBdJx+oPRBgvp+xdYGgMxGLrnDWLJKz2wHV4Nbwsn2GyRq0xJvMddNtq
+BN9Up92Zed13Wus53sUnNJaDBfpINJ39W8/Fb+YL319S6TUZ+eIv2wbzsvm9EeQ
34ddJxkI/8AZ4u9aEgsyBhn80/BOd9idWxfoWtjYOAO/d2/d9IXT3nY9yqDa5Z1r
ixDvrkwwp/pjXqwXG6NDOv7sxoEoUUnJr0JpIZPbpwdvomM3MxZNLo7+nabX/MKf
Q97Kkrj1NzhzifGtDm4wPinUmd5El39TYup5eznnL2tRTb3lhYVUSO8TPdCpWY7u
dlgoHx04nFPpC12U/DLdpkG9Kl4YfOmQdCM92RYMIKHfZADT6cicMDeleGdXkuba
d4GJn1pJy7bdm0JHNQRW25WpfdY2DnOWoxBzYuJBy8O6ZJbawahS3ZONoPomSgx5
1uBu3k/uhapKQBGWIKpEDQfMaTPS5+oDevZIX7eWXSI5W8A+uXW4xUZu7WVPtls+
xDxnlhv+oTaEr75zSaap9lPBedgxe0/yipaiDBuYCJVW3X90qx7IgK1711PP0liN
cW68oFM3VD4CKFzUYxEosxASszbMlfVCpBLhMZoBRyt5tALo6bUDa9DjJUN5S7s/
UYgI1NT1F+OT4+A7/HKmLWm+Wk1HoqGqDeOsjVA9e2BfdkI8oLt8gKl3euwYqc+i
lCioR1VRR01TG3godKfEvYusKiDJUujAUC+f6lzaploIDjmX3c7ZXNnF7VpR7WOP
t/Dc68YuLoxOsQrnbMOAVgaE7Ni+kcrvBWxBuLtztwKMOb33QMKR56VPsL8aPp7c
KBO8lv0joLRrwwlT/Q9pLjMud9EPOrvm5lHnzAa/4FBft3DxKi1bRd5+TNgawqbL
CIGVKK5LLio6RJNyV4WLrNWlxzwOaxOimQG1hr+zvcyL9eOy3Yl94ffhnM+xgd2v
nXhb5axBzMkvaKUJhIUoEWOA96QNO4RNDb3kaju3dA9FFc95djXDdsx0y1XcvkWx
4x49NkBGKO8VAyhmDtFR+GwkQJU6SXaqRDhOy5aPIaxTkJ3uPRFz9q5zVG+u0QUg
8zVjXoCBM0Dg+ZWqlBr98KRRopJ81jskhN13As08zTRE6rY/TKaTlA3eNh65YBXs
UqbnRalzkgiY2v8QCH5iR9OskUUmAhUuok5JmRjcq5k6vyXLs5WK+sd5JWSjVI3z
s2NN8Qgdw0iGF8D5ZS+QsE4A3IaYOCPx1hZ+2VFsXT57YqNQDM4k6UwE1U1lgohK
Q4ar4EtQ8oCfsUx6WRXV5iUg4gRW9wYYWG216SrGVqd7iWHiLlqcGmOjBtdMmuXx
ID7lY3iT1itpZq4iUZuQI3VUevW6nYuPBC7URL3K8+J9wRe/VLANV+GfshvtdU3N
DnrkcVh5pFVoHd7nhMHuyUTk8903Sz0yebijRt63TQ2hI6ilTnuMb/mkZ+t1+K/x
hmKlh+2uuTSKMTexcDN5BEyVwAOXvghyXQWoNNmIBvWBNVTlNUF3QZTzBL9L2KN1
ybkIhKhmEEb01lFHgpbXw+gsAUMSMkEJc9CJe/Kcb/Lct6xUj0XnbIueISKQXSJC
P4vM1WFhzyWK8Qae71VyzscmEyVpCglJn7Db0cD3p0761oh75JJHZ0LImp9ESpLf
7kTZnYC7nZYXu1yvEKionzAh5gx/CZYy6oGGyw2vdbAPjbPeflaMcLM6GJEn13R6
OoEa8DKW1RfhcywTvnMecu4vkBYdl7pPyJZVawW/3QeBF6lYN9Lfn97t8rJRRbsW
p1WABdhY2rW7WJUEjQyq6yJXIVxj4Pgnh7SQT9gCnPjpqb8MAs8o5jl8y56si9BC
bg2PceGCG8TLL1oEaEOOw7V3Cs2d/iekQXCb1wxYP5GvgnHURNZ4AF58MKlzLvNx
0FJggVbSR1m8gCZT7SV4SgQL1kgwUdb233X1DxkbtNyZQFYZDmbcrpna8vABtNDa
W4lSZXG+HeNWUycNJ3h/cxLbyP3SESyw/n3hyATV9ACtH+HCrOsFode9QdmCTMfH
Wy9RucKnOmBqUlgWPfxIBUtejuxl98/lRSe47MtoKA4RbZ6yeXQysx5fZfhvdeOU
zGwZ0TEN5n6KF98Yu5yWZxXYOifU4gdm7kwcqqJVg02PLJdgs50/BDQaZCFHjbJr
1XQGhLz8egb81NfdInbcQrxiutswk8HMSZWo0rdPPQ4Wkr0+NcioPqKu8vUuMm/m
Q6YfiyEA+RPV1Re3P+HhVFfhxtjpojmOar8rIEJmRC1RbusYMY7p1dQXGOGVCrXr
QpDemChza/ffmcV5uVCIOEA3qAbbI2apJNfY37+J3kK8dZwuC+Jg7ZQFtQteLSXW
+/JywxBcmKIO80JV9J1HuAv2puRKXLNlTb2VGpGRgJMQ/WDctg/YZJHQu/nAbflt
fBQQY/vAmpF+RlgOkHM89TC3gDMDraWgsv4Nrwedx9MR+Sdd0Oy2wE8DkZhL2Hpw
8DNmHzVQVgPt4EYcJs+Krab+y16cj3bIxTONtO5S8FoLjrlXbu2PiewD7Ua/T7m6
0w6HI7OSNvAW3ZRKUoDsaeSttW0iVrUyl4J0wlv1wvJ6yq/hI2MRHBpUZ6SuqjbK
H2bk5smta4qL2LY8m1g7deUunF/PwJ1QxpXfRCsqm5NIL3zFyetWU8H1PUK49/36
P4K/HJ+14lBG710elldzkfFQ6WUeQ+e2FSBvc8XabZZL6257xP85/nQ0nkd+6w+G
4zSjdJukd2pMmwD7HY2otPMc1Eg2yvpz8CXjlKerSSsBg/8klow2bMChyreISfGl
BkCxqT70YFiAAxgp2t6lhsAnuDGbf4blVnO4V4uzjx/cYyJumko904vFFS443jsL
RDl7Pp/JuddfUHKiSVObfD5QxMc938agCGkiUewm2snCiJ7EfyoMmUeOwTB5Mbw9
Xa2o5Jw6+51ePziec+i5PkNFz4FeIqNKlLldZtWfAA9z3ZiOY9H0RBVj0Sj1ogFi
wpjt4LIpDvopmXnYUpGLcAixCJ6aCX2JsRcbERhnJN01SB+GzpK5N7fpNDg6+xwr
x1nPsPfCVjE4ghzLmfo1vmid+9QkgFtAkAS5EjkplEWUGwmdGdqFD0QkyGskPonG
wio+s6MQe6ywJBzvpx1nBzfiLioMC/PnzV8K34ZOokBOtNy0zRB4giBtC5YyzN6U
Y30+6+ZiPvA87R/Bi8RkIqTVzGsI+w0hmUjaIHMiE3CT3Aert55wvx33xG1XCZ28
MGcIPIIBe6pynPYidUmaoIYE8H7K6O5oXLDaU3v05WRWXR6CmjSiHUa5xFnTUed1
0irTbuLptCnBVs1swLIuDfNrUgxXB1sXAdiez9LT0NZhi7si7jWWBD7n7Vc6pzfY
hM3/eYkRXIW7b+FbKZjHhLu7Q1GTY5kvPQAAlWKpT2jPp3BlDCvg357HZKZMauF7
OhCPz4RgON82XzUA0qc1cfS/WKUi2rrEVk1imsCiJenPHghxaajZ8ogfOg8Rg0Wv
yfdjaXxpVkNEKzOIe3CMYQfD275+PAcw0GCxRTZqikpU8OHjpPMRJ1YKHjMuYYRH
vHwkuO9xOM3422VAHec3CsruwFboIQkgj+sEoX3XBMnEIhb27Tm7FBdyXS8lmBqn
e+WH5Czogkmi9hhu2SpEwz2Z5yxQ8+OmlXc5gBDxwsaJebNJhztzyQmiKldUcJLU
fPj6JGDxTvqNsLhbHBVl9qonySEAjBnbZs2ifqnr6LXHXOpI+78rlYTxWIM0ARJK
BrnebKTKAk9S4SyFdtWVUtz+aLM4NtLwNNN/qfQVsjFotvM7FmrTs3FMmBLnhiFY
uISbc5g/Z1M94C5yV3SGRHr2BqAvpB4jMUJExys9ogK495bZOQRyG20Z9hbXUPUo
CxKPhfvh1fJI8j57DEmuY3xjIFAHtY/NIbmDBcoXomStgIihJh66sTYFstnNASgb
ZmKY0QBnaA26k/NZZFwvhyTyJ4p2SerPGWuwpNQI4zJOmR6PSygLjn6ReiFD6NE8
0haIjKJaAgw2a311dQkEGdh4kAyW/gTGDCDP/16NBlRvHpqd0UnM44S2yoPQxM8C
zhRfJ3yBnHRual32NBs5l0VsfkMc7TeQvTD9SWaHQ4MxAFBhcj/pItHapMPURG/0
Az4iXIBzk0lW5mZdZIclvssggKuThpK07As/fmQ/FMZXuvhD1wxT3zjzkuLAA/nL
jRu2BLhV3g0A7ARaahBv9DNG3CKzxMD4RWwuPs8G/j74IJT5cXo3kH/Rzt5vkZ9I
+xuvM8GfYO/f735EEfxG2r6zFTB6Pz9y2123r2fn8+fLFW4u7ZrWu5p4BieUnghq
AhwRUfoew+y32HU0bOFDaJukSollRqZN2UjUQ8ZqJr3Vg5XLAq0DTpYBkBN18uzI
hbTR+l6DLoGi3L+2SmE/yYUKIrYkeKUS/HrGI6qhqE5LYj3cYoq0IMlzr7A+7aCG
G9hl+aG4DEBep6dUyAbCC/U7i/1Jz8x299Sj3pSMk/Ch/GsxegGm3anjJToEd0uz
Jq8drUUJzSAB0GlPC9HgueE5RcLs7BGLHIwSoALjP5iMlLsM0YEH6hV7V3o3XCuP
CShjopsAuJH7jJ0lwRMa2n2Kt9UIYmggWBzhhQrNTcH1AzimhufA3X/Quh0gUO2S
l+OJnY5T/paneI4mcffHYUU+j14mNe6oAKAuUcmpRYXBqMGyO7SOTwW97oDRpqpv
HqObi0HBGcgl3Rn6iu8VV5km6qtWxuG6Sy1pDiecH2VgJZhCot0T0FV/FFGGMC0Q
DjedSIpu4FXGQgZ4joxnieXmEV6dJgB6QL6K+PyEqGGODW/H0lwvas3Z5tsHe+Cc
YmPxda4DiCGJdXuZP69uTXaMgpU2kEGoOsMMX2M7gHiYwdhkoPV0upU5YUjcQBHR
Cl33rSHRCq19ao21d2G17Z1ZZm0MMRAdRppj/TktgatuyGQXclGVb6CMDeH+6c0w
8hUnh63o4ldN6UmwrYlNB5y7pmHrlXgsV2UvEtQdC1VlCimrNGzUe7SsyFWeTApj
2okAo5UAzNcMdz/xsyuutg+bvHeDypItCSxLBOTLBisNqaxxN72FuJ3ChxnY2jeJ
7mdaQ5hIsqthLigPTPhO742BwWc+Ggg2eUFCzGhXidQeu/TIGhlh/+N0kPgylJal
y0Cu0s9TgF496CRpUUHRP5zBz/PtAyw7tIdPsDSDs2Lfpolrg5gkRglu+MXeaDGb
R8G21a0MpBB47xxEo9ty/koOe4Ud2zZiW4JIwpoJdInqFXQGPVVsM1R4U3LxKf6c
DrvkDNtpW+B1I4zUWLWWbP9JlbPNpZUCgOFTVfusMCnLccdqGmZ5CSN1PfpzqXzu
8rrBzSMmONe9oWlu092X8OJ/QoiUWmS6fFaqVrxQKk7QQ5r3JDiEcsH2lah92OV7
DQDQE9Tg7wRGLloKdj6hHr2bm5kmw97TkXa8+MD/3RwlBcb2nSXktPVsqsW8/2uf
uJB+QyyrhqtLIWct4iZzv0/FAb7Vc3tqV7b3kt9n6AhZ491gqoc+LT2K+po/gF1u
p3HpC62yLmfH4Vz7T2/fuw4FLdN8ceBVHf4A8/ZvBguA3kpYjvHWW8ohqI8BbuFg
f+4LwtA0Ys0tHxCUitK1geeK7y0tXzfXYDy+UPiVFb1E/WPdlb7WWfXTM3ghAAJz
6T6UFFVrFYMi50RKv+UUJF/8R3EnzPY2ZaOoDqAHRESQB6FwiQPhmgejo6Wbxbod
TqRU0Wski9Kyd96V2NC+fJ3xkEY1uO7mP8vdEQs2hWB1bZEIsaE4vsy2C6HJoxYt
9JWhICdV3uxh+23A5v2slm2sG7Cgw7omsOy3edN0wUstPSDEKQSMTWuVsfNS9NOf
7sVFdH2Z3c7lrvMR+ZbLbO5NAsulhDraBxpylgmvzjPtiIOm+zjA2KKYmahtz9MG
BLIercYmBZ5wgxW5TxNhapZdFNoeNV3ABiHPQD0pwOrKWGvEQOE9usc0vgQ5FjG8
hsKS6SO3zPyaMFXcX6KJAcDakJzQ3ibmSIcWfimcdFLkY+fkwjJ9ukZqZbmxBviA
V6xrlvCPyH2NS2koVe0uaruRN8LoDQsNUuqo9BvooEgnmXPZE+A0jP/CuKRlpaHq
Ao9CUwEsEUsCrR5qR3ioelM/tNTreC1h6QJqJPdVUn2Xr27S8xPJKPS9hHIvpJB0
yUzqqaQRNJl+5QNwJ2c6lAlhNAOFh4PBarATsZOuZTlnAOflQyNDbF5ef+wBCx8o
dG9GcU/qYszC4ogWkczZzdryxtkxUgqONZByv8WcwtaMkIqoh9BHjPjRjjWMfBca
aF63cUKTYCv4TcvDf3iPMGG8CCbmAzDwfUL814ZAUbHvtDxVec3Uyto96nD37Pel
1ElpSzcv/WF/pKnk4t7Itl6mhuaHHEl1A45zr9s4eh1KyLrP7jquDpvYjIlzIRpb
60KEnhhcRXfBAO/kJP2YIFkE/AxPGx/HkWD5z8O6fP8TwazUnX7Qa3e746EgU8N6
2tceD0POJMRa0TDUgWTWLIfzZXlQHAMNZ7Sg+AuPj1YaMd6Aw7sN9ovtVVIskVdv
PainzocsWdWq0GcuSwXndk8557iSeaYNeF/Z1AczCwtgzn1N8y5sHsi5qUtqy/gS
+JNJlnuYg2i1kts4dGfmkydLFeYumKTMLi8qAI7CMomZqfeZX2sdZTRipXn8k2qb
LqNjNU9YEN7qO2iFCcTCEFI+mVSggRhXwDcUhBflgNSZ2bGSxzHpisDr7IwkzraW
OC7q3823H6N1W1Gog0ECTp+g6TuK70GYUt3Y8wOyqQzZK1ex/jIAhDsmChpZ9muG
9/SU184ZmlyN8djNwNlneHbD9vr/GWMlvZSgIGSpWcY57KB7tpPiAQolzC/xEF4h
EhzJpPHKn8jWj0RTV6w31+HcM5E8T/UadN6wfvGEpHyqlFh2ekJ9+pMjI3KbHRAp
dZcjhpZjWxEck9EQVhYNq3Buf+6WNqUMkN8J3EuRyQW81RKYOBG1vLJFZWp/r7uL
7ZeA3vuigK+WMu4a4fCMc6/SbUQLm0Nj6D4YRzfgpV/KtVBLwoKkqCeQEgJbqxDe
RXaXaqQayJeTLKzZwCw8mOKbmjYir6XuArrp+iJoniLlcYWUTamqJ4qVKgviZvjk
neKb1YtvhZwUQGdHwdUWED/4jBYnQf7Yem0VF7h2BckA34z03+Zd2LFP3mA+rbH5
1Q6J1Ap4W4kV+K8zVnHC1qNkN9O7lbUsxUXcVjD+/KFzkHwsxu1Dg+qVDCeaR4VE
UzfpDUYaaCObtmqLpcKqjEf5WdAne0UpZDTA/GGURNZBX2/hrPifcPq9yVR42OGN
hgYS/yF0D6QoSIoemXNFaOppV+WDigMpkJNcwMjMKJBXy/UL5IUSLAadKbD6p4mQ
I+K/TVb4bSZd0q9RXlxfpX/yGWgNfL2sq0Gl3oSp4UzpqPQCFQwdd39LIRzzmXy7
xeHqgR3tAGz8hiwvsvjoBoHwQg1C2WvtqBn84ESOjRJMkHcGZLG10MwydjYnS0ph
TO6PJGhxhEjCX9FlRo6eU0r8GJq0dELs2TZT8uS1gDKALHkujw6hQklTlXwGDthJ
I4t3Zr7zcuhXqHLmFqtDEynbqMe1yjzzkhJhBbh7A2AMq7A5Odu7NBkTcf87NsUP
hgOEr5TY1TPjXmFG+zkAlrGHemxathp34M8mpw65PlZ//7aePiU0Q4HCcHll8Pg0
J0mYIcy2S3JMim/nEtkD4Ntg98F2BAkQMTWlMxQMnP3DmieZPFiQAtG3Q82YX39l
msDnACyUQ2F3BpD0bcR67iuiwDdiufhhlGqQJ1nYgdFQd0eGpEEcNygycykyClv0
NEVlqtT3Moe091bAvcJSx9FXL1F2VTGdaXZ5dZLipxw8MIQYakglmiQeDCCKlW/L
lW+1o/zucPxb9f+J32Sbw4YMHsAHlahhtr5FiHS3DMfpNjRQ3u3DQJ1WJ0xopdhU
UPFfJy9vMbyzv5HU9sFtwhAGvzmNjvc5hWnUa2gGasNGfk8jtV4XyB3d2r7RirR1
7Xcf1G4GlsP2Gyw9HM5AQqyy6KKePrWVLzKTQ12rddq5eXTxaMiwPgIyVrl4XMnH
ToeUq5CW69uH9Bchz04iJ/PD9msCsgNbXLVKJgnh8polwbVHZPIRLqz6vEKd3vPD
lQTUjEPfgZzmylWnkOKyuv/DMaNSNLQ9M6dGyfv5vxiALK4wSy/raMrNks0SequB
fohfdUxrt2nnwZPuHD7gOlm0UKpCUxLZ2bAvRLy80yoLBkQbv7LCkg6Bi8DbQ7Fg
QpIzxYRhsmWu1D6LTsVPutqnxpj8LXB86NJAu1SD7ReeYTceO5bwYo4trt+VdXhB
1KfbK9AxXNU5nk/9Hn4tLikEbdw9Rf1hMtO/hVLN4sncmnPrjD4KB39zi7wyfdAF
VaZckY9BunNAjqMtS9sKn8qvr8NHFzP8L9na6d9AxWsvJN8XENteoQZZEMFTZLSg
ThjfeNtdvsh9sJ3zTDnIGA6yyZzmfN5KF5vekbiaWew8YX+HdPPohAZBMHLrqRwR
W2cPK1RJT4HH0L6BGN2QWZPBO6C41U4m6P7gWmCYeSPsQBUtPmTJ0/yT+K8EqHrz
uDdi95uADTgXqGZDR+xU1t5ZwcWRi5nnl4GqHAJiNMVMvjr1r0nZM+USH2RPm9S3
sGvlY+C5kgYxP1MKeU9//wbvYks1x3lGIdU6TcfGEB9hQCVM0nlQwdpjSvuJGe2R
OwJ773VBTcsejedobmj/+JtZKEPCxqXOm5jv4FpjN0ovCSF1+otGYTze5vmh7kCJ
d+ZZsBybbSANT8DSYdvrB0xWJ3ikeA9XTVEMeADWvIvLt0LZLqKGZUw0QyAdHKni
YXGWLGnYiYSPcHvy8FEvM70qbrPue0KQlid0S2kMzg09m5E8X1oK5RF09/ZarrTV
rsEwNe1fwYeo9XFLwFwa00AEJRena5zboFHesoFxx+Uy21utiYS7Y38bi0blnHBO
qpW03KfTzAIQ5zDjB3o5/UemoTZ7HkjEFTQuwPNd5mBcC00ZYHE/eltNuxr46+Wo
7p99HAIxdvXn18evsfNIi+E1E0rtjTQ6Eyd50AP2Oftdi5yaDMQ1FAxHKPhlTkI9
Tjtq8QnvYPMNzFLDVoD2a2qFpPaRfL5q7ivK4i0E3ZM7aUahUwtwunq1MvyPMcUH
fbUIJ4APG08jBh4BOGbGJJrCk2EIOzYUhszQ+EegKaIOkp0NElX+cGOhTiuWveyg
a4sctQgfL59nsos2HCWT+pWCtP8AglDtvm/tkHobfFb/rHkBYgnBwfwn8VGiRxfE
e11kN8PuK17gdgG7+1v4N7s7OwLcbkOvmVBZN9c87yFFZNYdpJJM3XNnVlAQMq/c
CaiBa+kz21Hx4aVG9mXWgBsk5ajcTWlYM51e2W1z0XlnD/QpvLQUGiSLoKFlD3O7
wiEPLwC8Pt10VB/brR5A21zOX5rb6nPx1nJ72y09Pzc+T5FgBmJZ4NGLqjLPBze7
d5WCjXHSSbpRE8Uv1YAD4Bx6WxoDHWm8QiCS4P8W7y9tYd1fD2PHWGltQdGVGWrw
tUWGo84lKqash9CcDfppdZ9BhjMUIQgylSBJNYzznjSA6rdCN9fIuJBxABpnHaWF
D/bJTEk9vHx1NrfEFFvmSC0gJDfZVCjbW/Iw2Eg4C3oszNVw7JfJPV7zOW9db1Dx
UGatHSgwMDyhatJsZdcXoeoURLSkS1CAqGiUUfsm9fq+NsqMDMYIj4LpdMIJRFd5
xPmLBIDryY+2d8MR+X3Mk0+FaQ9BG1TcVUt7zAcdc/SGgKv7nYdHa7mYFXN7wAv1
GH9qtB8w/MMvFKVz3gXqZE1BxZt+qte92861x8QQ141nBDtjwTUuabPfSnkB8Rs8
YjaxAmhBHF480mksb8/vWYV79tJS+BBF1SUUQzlZwPZ1LdVY6OqQPPGxNTkFTX0j
j2j4IRb/H2QbpBvrVZig0lre+vvLDN8ctieA78RjnGmwY7qR6vmokrTSLvtuln+U
ddAJDC4pqMVOaN7Hr7t7Y7nCH8gmU+V5+SR0AN7e87reaO9PghviwJnzUY2HWyn0
7WqavRif43XBk3jF42wXHZzTvUsET2+zM08BO5Zxo1uuif637ZrIGGh1vBBsn6yP
4WhWx7SXT/Nn3uwOjtkh4N9JI9OxeFIi4Lsp5tuxsVb0bCcFUhSL0SZ6uw1/eGpm
+zIToL3+ju2xKYfQ92wA9pS3F+X0lgMdByLjV7rm2kPrRWVqzCEeupkDXiZDtiZE
g4HZN0f41eIZ+2Gra45rzYG9j3Gif061PZZq12JmisHkfPXcPxzZXcFeOvdRtDDT
Y6tqDqtD7mEzfXffBOd6C8ilv1aUh1+0vHpleT2o4wLwD//DL8AjU/s7hsCsjsFR
kh2Mwp1Gc5ifcaLv8ZH/fH+Wk3pIBwBcxiUKoOQQ7BE9F1CBjf/wvyqipqDa+dUf
6SAn0+NrIzeBcZxvN980RdMz0DUvxgknnS/+/tKgSrGRuq4tDvRPhIyLxAOr6Jnl
HYoXeUXPShugovNotsyQntpbVOIU3ouSD/ATha1eRjHEq8d//8gjbkiSb09LYInO
zWNUlv26l7UbCGjt6dCrU2fOLW6/T+8uDmTLHIRrHH3i8l3KZm26xQonq7Ms4Yo1
kDqrL3WIkmXUsoFmJCMTYvVm/O+gRKduNCnOjnqkMaXoDaT6GO9FOc7KyrimWiQ1
r6Y3t0mTteKTv+0MNoUGqJb2V0eN3r6MmmToz7mvpTepv5w8M40KfW0TiSxb5pXS
onUexKturyDJSo2itQtKXjcuFT6noGo7+8bxxiME8Q6m2M3MeCLzceSnEN7DpSv+
C5M9GJxGWXRixqNDeH3Hyld6bso3osWHUXU4foR7l4o3uTwS0Toq1x0CUu5JhHum
0l+sAVHImyR3ct6J+noxtbectBtGAa90ji6e2kZyItzKB2mi+Fk49wxskTiMK4lK
wtz1JzKzUKh3jS6wP2VXs/FBALEGEA/thWSKWRq1HILjX507CvTj/bnvc+PpfghF
9BKqh5ZnDIj3MaKm1mmj/bfeISyrma33UHpRvrSqs4jjEHdVmtkth/ntfoVmRfyi
7JYwqjACpIMcAUyVmug5t0jvm+fbT1ZriWIqjx25ywZYe4V0zkciYEHYYZWSUJZ2
ycJQ3zLlSNUnb1wksmJkUP1bB5TheZ3CZOJv6DfyJh95B2O8NkfK6pKgqZ7bV6QU
KlXhojb3is2GXwnJkiCpIN2tkoTi4KXPVJbXBJDTaDRDLcoyNdh2JPFZZvAWHz5T
0ezHEyysfumAyyQk6kGZIKc6wnbot/ufQqkbAhuTS+xFNctZq0TfKaQzAX07nnyG
5DqrX91n7P9coFFKA+jHXWavDFIrvjPGEFrBfz56Bb8M0zp95LtQ9wW6NsooCoYa
9yAga3frcFgpKp/fDUX5FYjuLFXUWzCWb4HUM7rl5lwv3vWL+pOWFtvpGf15i+WZ
ZtS9FnV6y/K9mh4R45ATc4W+D/E/QyDRV+VGan4YrdUygwlH0Df+NsJn+PlLWOKn
Y9fJZj0nTrOG+qepXvXCoqJjINIza1nKEsbv+MEPhzdSkSA7ixaa05gYZG3Mzdlc
RWRXBnKXk+ljvHCm5eoNWH2BT7Qml8SHaqpscsD7PSveMvtnHIL7UmTRsCmvHFcK
mvrmXBT39GNZpzJ+KG9/ZTqKgms820mDWsyamIRcRn08L1eayD/oO4azJOQZ4Vyi
SrvGb/A2wWoqcP+FUDzFFSbpPsFBW+wFJiZwbExBl81cv7F0bycfaL6Q3uM3kjKO
qetU2JA5UKvIM1iELqZpb0IJ0pZIPZWwBDZaAVnCxkTXdN5RTc9CLO5DAGwz6eAg
xofUMKvwxtEa6CNv87XlSpLQ54LBwt2vxg+zPytfeTx1PYlnUv0cjqIAIZbqhklQ
PFVPbXt4+zVLRSxQgj5jlsFtb+27hJFinCbExz1vamxgij85YXpouis57cH8paPy
fbBqYsw4w5QB4mKbWh3LfztCrGjbKKRD0XyJVLdpupxj//mwmpyo1ZZYTJSO68sl
NQ5clYSU12b8IWLf/S6DXdWQC68ehR7ORv+huqw8FQHuOQsfKXBtfGrHgIvlEZ1m
XQ4rO4Azx8QduJBDcdulwdNMZSbCW39tncPg8A/a+lMM6CbTKIh/ASbNdGiR1kEJ
HJTfaBz41QL4rgSS3zm0Ux9lVN9d44lCGyQlyQKA+zXkbXnup9D4XMu7jOQOjWCv
xTwBDQ/aNi1vx2LKj17Arn2GFYaZ8gR77I/JOj/4oLENzw4Pz4ZJGGpa2oeXUBV3
roqm5gXOfO6zLKQogoLdz7LnQlezMVlvBtq8tyAWsfEtQ4aO9xOr83gWVMjXrdOb
5hfkmD7dw5Zr45f1LbXmmPFoXemZPgLQ46vNvYrTZAI1iR4SXzVnrkhHzJGwtSJh
EjqF7D1YzrfIf1fW4lVYNMHzDOO3pkn6vu/EJGbDHeOaR00QZxrrQeWJM6QF3mN3
Ow27y0ra8VsYcFE4wFlJElCfkzBXu/bQoE9osasyT1m98ROrFGC+LG4pHP3odhCk
zGUb5W9jkJ7UytuhxvHQgRYVgj4EvEv9llKlsZBOzsZTEeG6/ptxeuZ7y3OSWl00
+Qa4R96kF/Z0rpR1zEx7FP4RU2HLUV8Vsv4l+6Qhb+f3YqVL9ZvGHaEheBHzoF6d
H/8zJ1LpFqRoo+C/OWSwyC0VlSF+S6s3m9gGKHAK3shMUROkIZhchq0CtzHaGLBz
JslMSdBCGtI/qs9RX1X+dm/S54OrxcCG6Fb4yJvOo2VDbtf9phfjXNtdDxgbkx/W
WPawynn/YUd1O/b5fil76juBrAF7GKG84LzDgdZd/Vymo4gGvETiNDyT5ShY+jDG
YE+7BAEwwrpJCgSl8K7KsMlbg8bbidxoxS/DuN05ef3oMsMJH+roY/pv3MjJ+RGS
qHVce5UoOQPWhtGzY1av9JFUmqbjgKT6JLNpRTiScBAqw9PwE+i3S8VaKwvgNy/1
7b+7Pf0MCSBL56rpir+mq00azWKyR5AcTxa1gqH4xTiJDjvwAROYyqVJAAWjUJ4K
Hq7HZSTKdzThKmbsHcqFzg+XxB1uABpG6Gdifvw4B2LzK7ArrGe/EWW8z0J3SrQu
/cXWSItg/vyA8hEA+J3o2E0arlmZBXfRxLB4Tu3m3jaIZ/I9u5LZJ7CSFqxBDHOV
RTc7CExSeZaqYeUe4WS5RvaZ2lkOnjBlKV1VVYhaynI87vjpYHT03R+hHC+KpKon
ihWsoEyjy4WGKURDcloK9hh3nv/4qDMKrAcbP70OLHX0AkeLFbUfeCGILxTQJnnb
J9/NuUR3/LFJ2Iy/xZOt05J8h5X3ZCZJ/CkTS+VoOk26IsdtZCUkMjpxZavUSVLE
rbAsBQOqe6vTcMy56PBfAhHTtDDzwaqjE1z4w3VGDMR1cIGpyErRYvn0F0M8h70t
NY0tMHWrt6v3xnLMNt8tLlbkV6RBhcXSO9igCqX8GEwCkIn1b6FRqVmglSM7rugZ
JSkSSv/uq7ptPUzxW6+R5wuKESaaXGsmUo2bu6BaYOVbjmgPMMjl8ZyVkcU7lfd8
cC3XyaitMn2Xy13NEHdj7TVQJkXaN8uZx+WoByqiYslUnGtXNhMDH4H+fmudwRpj
jF6VQTyctH9n9I+Jrd+Ss4D6cMbtzxDKYpqIUsM/PLn5eWpRTundOeZvZxdDOOGj
FyIfKaqS2iILQBUmjB4nKyQE7XMIgEIKQdBFKGGWUUjUKBeQWXUobn9inogoqqB0
/wd20cmQcgn4YUIpdJQsBH2qxcHHjszOG0pe8zq0OyIR0Dj+sDp8eRHirNt+0JDT
/z6fJi6tOca3jAZ4SMD7maVyYQvQ7ETxQOiRuBualgcspbkbC4CeajhDh7kHc6sn
na5gVfCsyqfAQGC0mTxrlTAQmt2EzRX+EY9O40q8qyKdiDlaMlvbimpn5g9/dini
Q0MEvVlZisUE/OKptNeenuncdIKWrekpGQc0S9pPjQPDosgLZlPX+WvKPLaF96sf
q9VplAHIkGwqXvMHOWwt6W/VtX7cpA1zaiO/JjRig7a2/ShESzjBsjH8n7duKNQo
JA6FiWrEEdRbLQ2R7DrdhotnY1IS/dhRwGLEIpLb2Ncfl5wN2F3Izq8fIDLGTy9G
qFV48KXCMB7xSQlCJ3g49Qu+0K2XJp3191dsaghAIfyot9QuM6T4jAEA5/tX9Wel
kJgVInsCiB7chk0MMkKMZsnaZg7W+zE+wN6gIYaSJhS3O/3rykYypJYFxW6auiJx
jjLFNmAeBmPjG4C4VNyildb8BgPg/JfBE+fTFwBY5OHKXWd2b43Qd01MJGJ16zqK
mwWHiFMSw2aKKNbHrCWhknUOwye0CGI8lH5btZ+WGKO3vq2qWsVHdGZGcoXsztvX
QUTHytSUOkpVGuLTkAr7zLeTYYzSBIPTMADAX0JdhTMomsgvOTAoCXZWZjhSyoU8
8Han1JXR0tpjiuWwDR11AhzDWu49LQ4O4UivAUOwNsbOdB8hEGj0l8PNuM1mtDAf
bYZJFFvBNYjzjjEuNa/afEiBwX30C/GFwXffux8QnqLf8uJoUDpPCxTJtHu30OeT
mwFHomGA/uN3efwqmUguV2z1fTCLlxaSwRcKejh1zVycsrO0dh75Y7BrDnQ59kjm
fdHELFkgpATcjh3AlhxGs3qXomWhRdZmkbB5iLtIOt7Gdd6uaxeY/mZ08Z0FutBg
/Kb+HCehl7tMHt7X6Pr0KDsCZdC1kST7sFlcEM1t59BVjMJ0W0bso0YTIjaPLZUW
TOR69EnIc5zV/uXuSzl3eQQ1pImqD4NgJRmxEOF+DHhxSr3vHsXySI2ejfY0ONmM
NXl9YfFGz76xvKz79jAdLR8oOhrq8NbBXdKh7HxLHW1tSf8OGrm3YBu9/aZihfdQ
mPf90m/OJWF3nERQ009rQMiA7oCtLHZnOGxFs1Mez+B9M2aca3yFHwJAVYr2zzEl
Yw3JYtaQaIXX+JFR/89zln79ZoqFaNK1+EMp1BFfuFRwTQT6581lCZUCsogcn9TN
s4bCyvCWUgbwu4V0X5ZQIqNf9kNKIbZr1zIZ96nR/avamRUHYtjmuvW8cjQ9AD1N
xPBVaprzxjhYQ3jkFBx7lyuW5ZSViO1kfOPNeaMq5vYd/V3B8+2Zpl9q+9lpJi5a
0T7r8OmSv/CPXsy03T0hsxkhGUSpfoKEzs0qhJkRyU5HypmgENB5EUUDDrcFzV22
Pi1vJSOh1tfJO0xEGLT/MkIvXvzRnNhJ9pIGURDX3DuavHanssbshDxqRFWQ9JUz
xgoPGkdstFsencx6gsTN7zgaeMehI3O8zhlCDF6RzXNmqSJ8aXwum6bPcDVLCmRc
uF/lLhUE1Rhf0UR72hx2UD5tBEkChtA6/gYzEE3IswczbqIKnJta9f/nCiD1WMLk
gwVrkPQwYBDgyAgGBHshjhekxQogaX+3nPjreYyBsiVamOaNx6qK5dCIXkkFlkoe
DshKQvxMD4rEo+OyZWIiYI6Ym8OGK3faqhHORRG3Q9THA9AxVbeWPwRcDgHyBAj7
ufLy9k9lCvSTNEiQWPrwr7Ycdh0hrTEWeE4m73kgiMBhVsbXSuk4OLhvft7GJUS0
S63+h4lwbt7c7LiaCsterB/DQdo/jxdrOgz59O7HN7FlTdElvkHPh3FhFKZmTiwz
0agP8nbl2c8n7kryrIvd8zdm3GTYAsE7F7JMNZHtOrWeneoHT+9Q5lZfIpeMoCWh
Xm7mquOMXu189TDeH9FvFeX9zL1+TaoXtb8eQi2ZRIJDwoaeFQPKWIlwTAGsAIBH
SIJDy/Yu5y3lppARFMgV1uBQ0D3zivwXgTJKpcFlyvuAhv9ayorEmEoP+y0NTRwT
tb8QBZVgkVaaiEIVxpwG7MHuTqKjJw2ODx8QUtA0z8ZHcnGpJDBH7Oa1dATR2IbE
SqYZgYqJ6Fz21Q3CBX+mindWnxmAcUVwCtAF4HRXYHiMisjkilV7eTLqu8G8lHBU
XdQ6f9rrE+9RGbPOLvcFfYAZ0hoarzM2gM7pjepUPU9WrIRAnJGlLE7OYn79HJ6+
mUmt6JUDfnQKJXz5eeCNdPIjaUkeMWAeZ0el+LNlXfIBOsLVGXJwIRnWH3inAlQQ
HfXvrJALwo0fCaAEhCXUQylu/yg1/+YWjyRfe4pjUDjqYCYh5VUsMJakOaEpaz79
BbvHlQcl0zfr+NHWihCUrlz1WjbW1vP2PoVHg2BCpPo3Ve5y6/eDXhT57zSWIW30
z0Y6stFxpmTx0vlGd3kGuYtN2OZn7syMhrfe6dOHJRxEyN7sUGTNl5CrspTlMLAg
bKfLK4hg2VENedKHPSw7dIuBxvbUXC46CORI1DcqkX22T+dmM3SbDcckEVefy3Cq
kn1Dno5QXg52z4/nmQyXk4B9m0v19dT4RdN0FjF/4sConEFls53e401uprBBJ5Tn
cOhwbpmjl8+gAqRpPMYxxrAygH56WB4NVC3uqkEFW4oNhx/yKFkpZITQYSTgcaTy
viwEMbs8lUSAZ8lBCYebVp4gUUKMwvBA0vw/HX8YjnzRQ0Cu7XNSkLGG6lTk2ugU
IjEWwmpm7DP+jWys6335CCc5WPdjxRaaQaLtt5NNjblt+Oz0ZYxZGtb0KZsRm/R1
/EWPjVIU3oAJk+psoxmBNnRVixpeQT4enTyhLm3XT2hTdFVOfz0v9QQsJwa+e7A7
FVE5G5cVr31apDiVaDfsmG3ydtmGhbaOoy9M7Iwn2jZCy0XjPj4hIIB0buF2I0Mv
j+u8hMNKp4tH8eHxDHuAnkRMX1rYHouHVtZdFa9e44w7SdSHRLgdngfEEKfJW9G+
enOt9C+XHMaZcIZhRalFDq5XCOt202QSYTiRH3ga7nPgFgHWBJK1608zDtkg+fFh
G98ggygrifVzslRiWVpDTIl66xkJpyxyHLDOBk+lGBC99DKOLEkDtB4hGNmc9hjM
ohz9Ec+W4w5ELsM7gJGptdxN77T6LqSzXcmObbnnmxHqWNbwG97gkPVRm8tbtU22
K13HlLfmFgNutwD2iz0vvdkz0QOGGbuTj3oo7aafIaZVXYbW4K0NN+vkv5VRSe40
0VX/UuMf2ZwRmL34rPMn2mhEmgFUTH0AQawQVYl9R1H2Kj2Rkhqwphqo7dtiTY3t
v48YqsGU8/ueArYk0EgKUExAaM7fKms+Cz+2kF+jh+UifAL9ejlk9el7iEIDSGdC
GW9ZVIyvKTydHNWbssJ+G0d1b7IrJX4K2EkmJeMnQSU1kgKGyO5nQ7Eio/Hx8X+X
SpTPmRtxMDe4etva23QcU38GFP9HJ1L5imUh7zFs1ALhvW+WGaVi1ylEaJ2DFnwg
7gt6u5O8vbQT5dGTksB1AjXqIE07izkhzfDLpNxXMDC5sOuaDjaf2ggOWGPzbV1l
hBkfHgdHCu6KdxbgNVESj4uOHpPrmUer0XHpRp4njJyEFleX3AHcZ1528WdQOBBs
KIK+KcHKnWpTpk9uVoV1DTrsRq8T/kZBSwsAIbz+JMaSBLw+Q8fVmZF0ITg/Zwah
BvngW0p08rD30QDLZDPE+Au8WltBq5oI5eA0WNc/0RcgWgqREz86/PxcaPTU5XhX
AULpMSLokBXZb6lj8gQ/78/SsPYQe2foj2VVPKKc1naORvv+TNDc852LbN+GjTwC
A00iaD3Iz81ms3KlQ23f4VBYG5HO3KikhBogMuWarDmZLg97moye0tpPGfd1oU+i
BeJAWPu1kn2v9MFzozvPrA0U8YGpjGp2rH5mB+gIXO2wWHcjoZZaTHnZSs1x/v4C
e22AbMNgLU3r5tSnvzYD3qHg2offyGCaYwS9HCqu4sbzh1bGZCZ6T1LMH6U7cRjV
6E8tPMLt/0xzd2c1SC6WA1EJUcsrnRUiNoAc5QZGZjZf4VpZDBHMAokCMKbJwrGn
GL5m9xrV6fny1XBIc8o4lkLMNPNkr+UW2VaPV0hDXQ+FgAaqKgVnRm0qyeRU3SlL
vQzH65NrrW/5H9HlGOLHah+5Av82wsXkPiVFltdalMqTj5z2Do7TY2mRWX4+mC9/
1/OZUkULNKWCdQQXFeApnBkLJ1qexGhwfmwY6TcgRlKUnnLEubEPHEh3huTKBqwT
agKBIAADk/exEhpUdi0Ry5fm8BWtj+7xZoBnCrCowIQICWBOiPxhFLGS331QFW7T
sOELMwMq/RTKm/xel1bVhKGdwhcc/CgDvUi6GN9idnJZvExVTdq71Sb4UIU/W4fb
AMX7QeDccxt9u8J3MfztF/02KagJglbM32v0bupVf+CVCSXBY/URNR/9zKsDZ+fw
Z0/6EMbN/amOMfY5jjHAcenU6uFZK92qiz7DK/qVUEN2v47FXRls66hV35ThDSw8
hm2WMevLF3LQuwcm2BqocM/c3NdTowdaw6BB7+ipjDqTk5HdBGv/f5iuoBxb2Uhx
RBcicXzrAAN9gW44D9lvjqxMm/GUXFFe4bTFg1mh0VqMHnda+WWzOH25i18gOair
AyuBBrKVNYLadSicOO5XbKE6G/kMdglLxBpxdrJPIIMXo3Q53NVsZkxxNxnvUIdz
cG4rcDSTdfJkph2DtBIsP8+FpIuQyEjntE0gRaEYlOKV3LDMiNeygUZcGPFx82es
fG9usB4CY+1plvqAUeAQ3ki31dsK5muKZjP32HZ2G/aj4IiJ3m6Af6CZ8RP3RvI6
5aM45pyctE6c35AXe3SmalxQV2/9Vz5jwvDYwDopR7wIzzv3fltd836iQD1FtwlK
sF1HBnZd89WApIOWz2FiIppyclleXAjsGTp+LlBUChHQWZdYKvA/vqs1Fadfpgpa
CyPH3uynVnYCzpyaflT57g2vLV3iCcQjls1zETA2ifgwOVM2nrnuHj1ECV8sUlMR
wMc/NpobVNdConvr462OF9YnbXroG0RaUT4g3J7Fn6gzd+0YwaGKXWmWK+yLQA3+
tjdAqN2PHV1eaTMMiCtJY5uN3URU+yUzJxABlCChJYFAQ5rp3Q+F4j9JNCBvUr7m
y4CitKg3NBuqrWzoVuJk/SAqsjps/bH6wnRMiqofTueEwc1l/mKMPvTAob6whEl4
bFsagGTv6JD3zz5QqGTJlOX0GtDwuJW/iFn9JPH8gtjziCLwXrWB5xQCXoHloxZ5
my26VRTnN0C78l9/K3a9vjlJ+Rlniz2ngCuM3lD8/mteiySXOJ8ZFgMlx450LOjY
skBOaiU4ODEwiyYvy6wudgSTvIN9/CHVPUAI7Xgnyz/tE+p/6XPdkKp4iZJGLSwk
K5/pZexYTA1oWeBxMD0C6/lfcGqofl/zCw1fwjQ3jdCn2IofNLOP03657Vgff/tn
DQ9CvDbgK4y0ReIlQp891Vi2c9w9ssMw9OVRwEBYMu+dNUwaNB0wdERC8R8adZFT
VL/tCV48zXlH67gzkBQW0hePlPSkc2u6wn/INUbfIQSrTWntnxlkBqd0ZyRj97LI
tsZxnqhZfZ5SONpmWWtZmdZXEYpljcBbw6dXwFJEVT46JftiKITwowXsUQlYe2K4
Omyxbz4YMtqdZwwTWwjXTuhzMahmA7o0dwcO7uvVlYTdhOFxwxly9N44I6N8pAgN
0Oy/iP325wL8zbjAuAaP9j+oTxhhpWZT0fVbk4NNcJCPsWOIej0Oj6R0CztK8AOQ
D8FG8pRr5Al5J8FaXL9JXvCq4NyiuTprvATTTxcck1yP1iBst76oCYBb+J+nIt1A
/TVom+7Evn0cWDErClRLohQmTCegeUOHvzCHPl9sqOBcH5Sy3fQzcMtwjqTNQBZ7
l3bqBDFrY6A3823V2ukEI16CXD72BoQUwmMZFbNz1e860S+BGxjhuMHorw+ihqCP
yEAe1zKTJSkLlWKTkjCN+QKezfufaBTiIPdpqIxEUHn+GeFPLP5XGC3AyjFeMqd4
WYdTirAsb8gzQWeBAZn/MxHcDbqb/dNX/aUicIVBv9YmOJTZQA2KIfsQLV7za+wq
eLFrVzRJ5LCFNx862iUADmFYrB2BI327j+hVCSeJTr+dQ6RnX/lg1/tTDiNoFZQR
hUeUXB2f9PdT6rRWzuwkYA5bhdpPZEJCcyFXAXqOYiPkzRA7mHuwc45R7ifMwfCW
XPdKQSK0RG1bRJQ67CUe3kfZrQJDvkRq8iMZv1wyp9sdx1gvjfK+CNUGjfU+dy6d
tNReoZQUQuZ3Dsv3+UYKWnMnKyqHKAEnrWStYGfl2IXHOVMKeYOfRKk/ooa7SNsK
WTsb3752t5dlTBSg8A3CH958KUIugtcqV1h8SaRPG5h1nEudNJYbsCWz753JgkgV
21qSr29XVYOWQXAWWYLwx3FBKDTISwSZCh2uJJ4zP9BlXmfT/bTxuHnk/xt5mGlL
wsLcm3lMcO5bCeKPY6jhdejm3p+TuclVQUrsTu86Pi9hFBp4hfGfYh5O6d2d1dDJ
/i0ihEBTChLM7kDDMIq/aNNX67JQvw+Umb+90oWV1qdtDBvRFkEHg5MBvSGQZxRU
pLZBz7NxknZKIFbkCGJndITQmG1SyKLukqwN9zVHi8PSYcwPQRRI8FC6/kLjpLNK
7S+Msb6fAwzP8776/FnvZ35RG+X7WvVd1T/gT2LonDZmdrE/urYzFe7eN/8m1Ndr
+C8IHLseJg/qILS+/296Yl9B/R7nLGvdFe1RYuJKL0GeuIkqLv6hW1bmGIEHv4zo
fkmE5sYZxO2Ic7pJcfh/V3UuT2O0UPK5HFdWhKe1wvgJABJtlaKn58d+SiEZ7Ftm
c5gVILI8z9XRwlbz1Lu21XupGE8DDXi/MtQbmISTM2s4726sH4SSNciSJu9dFLIK
BUzlJViOUoEGQwz598k9pNTD4kP47Y5o0kFje2N2hksadjv8z7h51lRhVGmpPDDi
9s/yfl1pkj5/c3oAQmy0y3sTq1L6ZqynjaXv0ttW5fJjPtSiKCwB/ocFoof13VWe
iT8P9KLOCiaSE9w8cduNa6/u2Kr53i+Fe8f8ElSk8gsUzsw5uz5GrB15UvtD2Cfs
H77Kzaf7afP4wqOSATtZeeEnS+A1pwsGVAatR7OII+82pOlDwJAa6i2hsPs4RWfr
i+JQd0fBpLpEJkKy9kpmue7aH6kbz74rDe0qhuZZJFNOvWpJaWWLQCUyaxP6QonU
IwaYYwUiUT9cGQMCeq14BQflkEg7797b19W38bnNdoLIq46zBgNqDDDizQLrHF3G
iLoDOQL1Pt6YF0tkiHCFehs7z2mLWaHSD55G+twp5Hlnx8bnO3lMPJaUfODFTgNY
dqlBOtsZ+an9FA0sa3XjdKglXdX/zgJbUDWRjJsY8A9nedHHTEjPbOtLw5yQAXfZ
ZO1ci79YUQyDlKDOcuw+7mEULu9bQojh/ANjAy0kcB6WPu5q4pD8O7gqUiJH1NWi
VPKgmgKuZl2vlLcToKakuz+uVtihqsDaFvqw02mqdItaJl6VV0vl7Tqy9vdsN6yd
1y3+Y/zKHlK1TxXZqhqxPxjvAMcn6mOcaDFKRpYOx/ol5Nuwmn4YwOIVGmU2T91I
XPuS6ITH+I3jIK+tGpAtQA8xXAmQRYR2S4PQzfIw3LAK0SesRBCdXpLzx47JnIQp
YXrFH6aL6OiMw7YhOEc4FvjS0JhoS/Y0qK+I3I2ik/FwiAquOBVWXLnXyzK7tAgn
e8Boa/WANPvo1pdVEJCeR0gao20ZGiswSa1HpUAL0TGmBFW439qz0epaqBQ6RddC
IOMtrHuwAwUbhTEA8Y1J+klYbNqCcBDI2TgTfT+3+gR11nAOUyvF2QLnDi4lWMz6
PF7f+QbR2sBOL7xxzp0Iesx1qtsdyV0HMaJ82sO29P2UWf5utngW3mAALpoIVw02
NuKILOHvWgdZyILOsU20CRDVulplO2ku3/Z8B6IOWypgKZMIMjWX3r52MCy5cGp8
feT95d8GhKD0vFymjaUM4YorG7LxhYSh3yEuI5YA8IXL4dJk015Qgt1csloykg8H
Eu4Me3xQt5fLyyBnNX8zCB0Yi+qDfJB8nP43/OG0F/vcihekJ8Va6U6Y9lPmG2R4
qTAPTN7vyZj3wymOUyaenDvvrnqTlLuL/qnB7K2LM0w9VsL0uohGYWKSdO9JtUMi
1vbrSY7/eAkKn0AGKkarSeTjoqmSXd7PGRPiyTlBUEGo4gZcZQVLxeTvVhkTwStZ
rDh7OSqeg0JFYnncONFl14GRTv5B6wS4qwEQzweytPluIuP+Ij71XvE4MDrY1rOY
FinY4IgaM79OghAj/bn4xavAeeWE2A6KY4ZcJXBXSF4gs6fqNX8JPzpaC5QN/GVG
gFm3ZySOFVL+q1yqtjGPjiJc+lrBqQOlXCHhzVPJZeVKZEKStAKyOw3ZNTzlHwxi
4/H5jpp8tU9Vr8UYrUV7QhUmXy8IshSvl1iYz8YsJ9q3IpPVhkSGs+wT/FJSa/fM
CjCmKfZmsT/9T3X4vTGqTxLFiQYFINq5HSFdb8/yqo6qNFQcEtMpxa17A/ioKF3e
pX+FgUvAdabAsLx6WiCQ9N5nfmM8HKkCS0Kpbg/hn0i0QYUvB6owGqLv61P95hSN
P6xsgomDZydr/xoQ1VB/FipGGq5Hb/F6quWL//1vBitEUCBvJOpIy3bivE46IqX0
vFLjMSdD1XruKZYZ2rDjvm2LNC9OT3qf+Ew2CKRtAVfVZOAWABWuJqUaSbOoY+5N
GhWlxMk6IuayMZCSh7fIC23bSePfR4RDdNlWSrGI0wAoc6jAZjdt/yczg6uDiF8F
FwE0mjRxS9cZTj9NzNJnJ9O4SFBFYjDXBhR8Mh4GhnH434Bme2xCkAEdtpWYRx8i
vETeEx4E0cd7Mf2g+h1KvuZc+DxTZ85IiNO4UYVcek5gJuJviNuscs6+jNhg7ERX
28NVbdX+SAOp1oHVc69vkh+S/1Gfldp46LgMAUS1syPN/9OWyeGgThPR5ZNdt8Ah
SPmT62As7NufSTVTZz2Os2ROAJ/E4w4zLljPlyb5xnNqTeBJnK/lUKGSMNxDqUlI
oBp2i1hg1l401mA7BlJVnP2R1esSh13HOSnM2kuGu2YyRZW9xr+NEk1uRneHtyrC
EhaX1p8PMLXJJNQ/5Z4KgumSmkxGVw0hllNQhAz9y2bLWP+3CuryCQqddQu0C1mz
eS64zO70I7J3jrIN1OFsy/DKgfT+42ANhHoGyUZSV0qdR72lBzuUxMRw/yKZjbCb
tKVa5lYRobCAHDsr82YqJN4hHhKQmU2DKd1XMGtcQoqEluC9rJKQoSpLT4XsPZA1
GDiRn5M4I7XNjPygBkDb+xIl29+W5zPaLls1n4+WEsXa6M8E0QIUP8X8Nsw8RpGX
vFcwBDR1jJaM6x8mFG5dumMJxaEirz4y0Az8H5w92xWaHWihiIVMjR3eAJsmMkhI
8x3VPYkGsuoHsVARqNvlBDumwbg5OvspDt4zua5C8kFr2WZPhyAPnStxUQbNZdEE
7246+XsPg+Xm0gF/G21qFf7wRi2F1OjRtUWGxa8GV1lwizMoLHhLQ4uJ293S9YVI
E78mNRszr9eHWG8HDlbsu28KNdmMA0uWzFY+v4TpsiAVBUvWhXxHN3zkGep9NrGe
ZLfF+hRAqO27FC7kRnZsa8w+7aDLRyAu4IdLJyPcP1WShDtWF/3V2klwtadKzOH9
XEPmYybUtqVPv+gWL2Dqoy8Xyz5RvMprOyKfokQfW0Mj4+mQGc3WBHiuYJmkpofN
vtAz1tTZL6+5INRqy+vcPEXpOQT9rF7JHhCT1gjNMkKvPW9IG5ACbHEHF/DpITC3
ULdNQRJ3l6tRFAkYuUrs39xJhs+YcEYsiNufB7qryLaIh8dK1CUR1+u0TwMM7Xa1
hEObLmlgHh9dc+TRN50gqzhL8dd9Yi2PjJfkJzQoGj+mp9IlzS9t/Hguo/qpc/Qo
5zt/0HL0wEoz68cMFNU7CZTZK9XYbf+BoUv6zbhg2cvLaUtykB1epO/yhI/bz9nR
zvtzuQAwM97vO8u2MG5mZSV2m29W1a2JrOsA3ux8Syr9fqDaDZ58/eZby7K5OCqZ
0KCE+H9yuY7iAfjZfFj3Tgikxl8f1GKVhbSjrgzCFoxp4sVvtrRxuOJDAe4JZB7n
V/YtDQr9dTcfkTSpS2c4hmExpGqwztO5L1FsRK8d0Kc0ESOc0XlMgBjKVY4/reHc
6ahL7Tjzk8cnp2ihAFO5uRhP7QYPo6sXtXjC0RNGfvehtuxBETLEzHTL15bfNm2c
8JT4WEB8WabQukW/zd5+lQJRUFPZy/HT21AHkAGx2jnTK3YC9mhO7gWs9dvu4vUN
Wvu+CbKYHLgdULoNHPVQ6V3qSTxT0pr7hF4hKd3Db9+ri35cf/ZyzPYzIC48LVkL
NvzC/4MD9DftSvV2YINBE2lmTlK/p6LpF60FA7DHFW0CIdU8QMHf2y0nmWeDLYhl
yoIBfcraENGdPYjM2LLNb4doxZIlaG24LdAI/BxPY+/ut4kNhAx0qq2xowQOEhvR
dI3zIj+2DP7enAKO/dp/0ewlRcMvv5D3Mfh8q3aq1ozCN0YA2X/MQfTk0SA1Jgu9
RFizSTdOuMmvFaYOjXgIDXbCqGuthuN5jxO2iuxUIl+EA/Z3U5PYiyMygWoN7FVg
kZDomDp4l3Pt3tT/+q0oihGWBfE+il2V4u5/PTUOKAfOyT8EZEog5AYnWaAIHRwb
QnLBINl6MF42htqn3pKcdyfsh4ORv+rHCPdivZFrR/UfiT5ayBOKtrguS9dCDFJ0
Ne3Tdct5+hXxKvKLUH0c76dO0D+HXsZlw3LpvjEcnMg17/0FAuivIjlei4k5BRTf
OJ60nssRLpj8sV6ZBWXvK6NsC2Xu4tKMJ8EQZQubB5EszrPRFgYlqinGT7dV0akH
P1vFzicOhQUnPyGMnXUSyHdug07RRRLF3ACZAKZjXfDHKqDndMLarxgELwnc6nJO
3Qz4vZmGqVEsIBzjEc4kglstTC2udRaMoQ8RXb7Y7jA0NkAd+noYszjHW7vWmuoX
0y7HVyrblWSJbvyhUc37iw7kvtCBWr2hQkLbYW2Z2CvfoGnYmhyjv91RTJ6Wlejl
4tAiHpiNLSjA8q7+oG2NUGzlKvNGMhHELh72J9Jy32j2yYTDL+Ttxq091o8HmIlm
8yxuqh8nISPF8KZRafQO+4bqnPH9CnW/bRuQi0IjIuLKUf/TJozrUMMf54BuIOmz
Hxzb/qGL2yXsbhpoAf1FnqVnzQ3Xlu0oVRXxuUk/5WmS2250McDrzysy0K9vdgmv
zjQUdASfn3FF2do6+bNVuX5F7RsDxo1ov3+EoF6vkG80IVh3b5jP+ejDAyIY9WIY
OBdpQp8v2/oxaI0pi0ReDU48vTsu53l5/Xx6oB+/sbk8dfH3BnqYC8MeuHtTM8aN
cuY1feuUyU3eoYym+nDzgLxXTExOQlxECLQK41KucbT4ACcotUk1YM+JyK+PFvkF
yngFbrF5+XV4od3eOTOaqh4Rb3Dguqh3Cq+s7s/FcixChTvpX/TN5fChB0ey5Vf4
+9i9UZ3qOvKn1+lYY5ViemXiRIFFAJYExi8Fg/8HEizJjLa86OuXG1sEn9ea1Zrm
qVEBOmt5Vniu2w8L/qQoZjLlPTSrYVNFup6Lgz11X2yPg2PiDt8TzXncVG9Q2YVK
IWZIkp3u2l6Y91dOb/SokLILos97QuuvWhU66lRYKwpQ6KxTQo75QoBg3pyHOo54
kWGlJl2ILlbiZa4xx9bwUCogDoHUXLLO3AgmMPqFgfB63uO3NcJEHZaY6A8KQhqk
lk5FcPFXoDPAUvnL0aiYMGfUAIp191I2OFINTKPs1UGELKDRWzyWgzjQed1ggLML
HTIXfL2j0ceNCaOvQuQJ590j5jg1ULkUAwSXpqoyP6mJZPHLde2kOfgY+CC3LtBN
otK9d3SCzz5aLu7U9vrhJ2ixDEN7848Mb3Kk67tT9pSYx0l+iWV7zl6iKxrSJfLd
Ih0AILabY1+B6AxGehoaG9Mih3rbj2zhgZJt6+bz7HDN14IBPVB6XyZu5VcE9pdR
Dg8dKjtyl42jqmq9vgKmjHYgpLNcoHFmzftSG6GiX59ga2Y4fPWuTJx+dCqQO5Hu
UfJ7awnclvc27WUvUOzPTx9dOmPxfrvDdLFIqR4CMoKovY9ixXSWTHK2vWFJrsH5
v7s2Ien0kF82MuW4g/dNzAzWLOkJl1oxfuUe30YyCQtWVtGDseusxHjTv7h+lrty
7zFrMnaLo73DAmu4JW5Q7X7mvyQiuhjkn516g/NjOto77pWk7rYlGNIjEteVt1dy
D69TdTck7b1g7i+8aR2JCF/C7ek1aQPJMK+k2RbwXkGLf8wN9+/a+QHJQtF8XOCl
SkKjTG0OkIQZcFO/zAq2ADgQmnzV0kDzvS9M38LTHxc84k5v++ohOes7Z7NTzxx5
7a7EeTSbfRK0WWW+p/SyHhs5mrBwF/GtN3MqhBJYJwL5v0q9TSaZjYrlJpwrKrje
h1qOu5r8YIPD4deyOscLfwSLUmO3Uu7c9EPUpY/L+eFO6hzd+DjR0sCnf3T3/vW0
/d0n8X/ECMB38rFIhjuVWlSBN4ypb6+u7yyDiDHrkJPxEENmtvAAHRdQsM7Fgbi6
5cEJUIjqh2cSgEUDR9I6Yii2BvXqx/nxXuALiiIYryGCqNPzwok9aWtYYvVVGwjX
sdS7BVzdYWcmsnyOE26yosuIPKoqLyhSjiMMuDUzPYJpAmgbNAOhFJgiI5IH1LAT
LZSlupPf/XhqDd+5AASJw0JGtF34BuZDTgV6cT+1Ah1ao2coplMp+TswhWQ4Yadb
cRDkHt7mdccvpXKJWBAfAg+pMxawIFDaVi6x9qREs7UwX3kst5TGZPvA7OqRgf72
QlK6kYHlKPeLKKRDAb+mwC9WF6x5xSYov6Ud++lmEBvcsPe0NkLK2LJ3OTXWymdL
36ovL66+c8ONiqMIq7UHt9xdGVS0cfsJzNQ29VxduAfgl2JJb7Bu2E35mCQ9FIKh
QK5nF2VGx+/AmCy5m42aZ2zndVBGuRlv3J0jOQk/uQY1Doy3yhz+B87woSLJYn/S
+O5hkh3Hp1FPU+eoXDhGIzccmFokXNUmlA4poDcs3J/kqYytMKncwRhtTIGwmJEv
ghz9YsLBTseVEzpnrGcA+R2PBSaSrU+A/UAZGQS4ZGbqOOFi6h6kmeWWYUy1+JvF
REFkq0/XO2g3KRrYNmNWlQdZSdzx7RCjqoCxsxKN2yP3Jc+8WXJNSusm/bmR99jP
+p5ghueeamZQuyIBqnctCQIHApkTp87yhcoO32MqJt3gNuUZ3NIgrabOMMQPeIFJ
18SBIc0eJX1p0bUP6RQCOxq/58E7lQm5JoWbePAQDQGQs+ACnwQO0ilQaf/IHVsi
DIjiVbIBMSsi7f/JuPas75nhjZJy319rwUo01Kf8QjHqVd4Md51SzikUEkBOR0kU
H7yRs2Og+rbfVNNoxtmI4T2qtCOzTJpr6a387Hmba7xu3thDahCcelD4WTyBlzEV
4m3quxgxUElxCimMWY7BCkixnCztHsQv9XtDMfUbrnfUneTj2JUY+2N6OSUHnS/O
bWab/7FvlHfGw4FHYhGUeSr6NRhdBlJeN7Xknn8hagn6Jz6J6MX+6EDtUrcqweoL
s9dj/ZWalncPtFBe24NqO4zkwLiMVXgrZwD6dyue89hncOhvJxZcVBpsWjmTAmjF
YpryaXjj0PdZyKoWhPSecumNn3m3Uh5645zkhr6vuCD0HjZNux0h6lQ6NWvFsuMU
JBM1+jPNYbVFiGwWTRwubj8DrD5i6fHNinHOSdbuTtLy1fISh4uOSXaLpURboWfK
fB9ZqH1fJPd3+afZa5z/FBDp9N2szb/aVQDSLSDkVklNmB8rpcZqu59EBk6bb7BB
5l7+SX6hay8pyTFXQE8eGZHTJQfx9pvmoJA+/H4f51NqD48oYBWjvSeLplvgessI
UOTuhcM8sPWaZpXJOPI0YAArHXeHmBA8/PqbcuvsqQscTnfRT5w2qJVM3QKFniCv
+VM9GhF1Fz51v6ecu24gW4jKQyvDAFi/gwxsMF58eScgN2Sf7LAOKcMoKfp8ptvZ
hjJbFor1Jag6ZBB3sK6RD0QN/iTLyhZ67RjuzNMUxSLS4YXnLwLxfehRGLrewzr/
dtyjMF+ZTKyggczF03SWFbDWeHmgealhITHLJpZQt/GH6GrwTtpz22DRjoRKB+w4
uL55VETuklcaL3+3S/eliCHRaD2IH1035nF9YzFqGTPDBrUCStd4kKUzQy4ZcKBL
GF0bUT19Qi4K6dKdRWKVRZB64EN8PhpBFbiRgqWhj8s8fIo7jYC6mT6fJzQ2P/AU
EipW+Ll8bhFcgm8PqdZinQyFzripeWLBBcfUNGdlKUdv+8evmezdvtzJiyz1Pz5C
eHV7Y2CjxvEjKLG+u2AFEAeTGbzZvLrxQz2H5nQGSElHdKrhQAgCfwsxJsoZTQEN
ahw3NK9PRGWI4L+YLQ09kQpeblShaVx6GhmUz4oDpSvup4WTxI+2qvruoJv8E573
rZClpSQRFtM1HVvhzm9eu+HbRiQwyKxDcZgS+xkmQFpRQF8S9ZnlRZp2BYeXBUzo
w47d/zM+2bPkN/JDLg0bHVSPPLAfm5+XRo9TT7RLguXwyDCQrj/Hy2jm2IjPY+hJ
UgbKB5X0f3S02d9ozgXaqkvgOdA93L2tpt6MqC6xLMTXlilbjZpRcX3gtBoIO2jw
bwH7+nUxhjaXiQ+NQ/0mjsst4u6KVgpFH8BCfRLGScwoUuCEZ5OYxRoQr3x7CHTn
stcGE32zw7NcukEXd8kzWisR1WQBLa1hy7e/Vh5T3Ipf2u4m7qDncEoUNdjCrlk6
6cO4i53SCTjTAp6KIcFDCviBPebgy3mQ0vEUv+RYqCo3CRZPX8BHOQXvMMp6LtCH
GMLZHQkszABnQRozhfb2EV7f5kCEgMthUja9T+989W+iuM6uHv6UgYz0yX2Ayuww
veruBmsJzeLIZfSAhE+cTfGnMuFFWR0O4JtXrBYPLdh9vGE1GwLC7Nf4T4GGsd31
4tbVJHggEEMrLmiG4+RoZ8CAnOA9WfvVFttIYMGlYrcz1l2oIxVdBjknAV7clCuH
4GD4e3rrpqQnUevEG4xD6+pibE954MfY9ZNMjwgloclntz7SvijBjpOeWo7Mmcqn
3GTPC/MLkQuUYzXgEsACPT4yvd14wz7v40WWl4FNFr5DJEdcv+Tz3XmEfyJyKnaD
7txTS+/+3pp/SXUGCRem4nq9YJtjUMaz7wOWYUQJZH8fdi1Artpg6XpsTjqBT6bt
NGFDXaXwYyDgt81Ph36ijZ7xpNT3h34Ttp8Tp6O/5/A4IHVlrSFw+mimqachrGek
7NuaRbVdxeKzBbZo0kXJpYnSKIvMB/yBqUc0bSKl/gd2vkjjk6UVde6JQy7dzETh
I8JQaLCKVinIu+eV6b7ics1i+0DByITeFbssIYaYbHl+O9SiQe41tQKyQpB6pwuF
u/55hgianEVp4sb9u1d+RllHHCi92TaSm+Vmxx090Ko9DMJr1Lqf9p8zF0Mcvkq+
wc8xwHxqJaxigRgWdKHwloZH7Y8lB6v8qCF2F5fA+4SAOkMRMiKFdxR2xdSNLtk8
XxpG5KHeJSbM2XplxZN+uui468gM3DPm/7M2B28GVf0KUsqSMr78zwNA1B/U6tKB
JoJvhkqj6YAa/vg77gvddw9DmDIlIuBRd5xpXI4pQcHXq6CbODuXyhNvpGTA3Ric
pNlGC0n8lpf2OhZgiUeg4p0Bt11PJKmZywAhM1ZjPfUJpQUE8BlndfhGqVrXCzMn
ah9ljR9J9PEWAYtCeLHDSKRqhqDZ+74Q5M9R3jXlGgzs45tenYct198MG8Nve6NQ
BSIgutWg8nindOl53ZCbq+jhnNqDsYFMH0qf1H4mwEoSzw+HNMMt3HmaONqdwSBv
wxEv1R4qt9LAsrFZOe9wp9P4vX8JQU29U5uptB6XNjrAMXaVsqEHUsuOigWvBGAw
V+6UQtBFHMhjvm2Pbwtek2HAof+zyPO8XQKugjZ2kQXRIMznNlZ85E6me69CuFw5
FJgaw6hgAuZs7Pm09vTp4GYZUd6UKM4E4V+KvpfR2cOGN9IbrbXYdgQWLZ7Z4pEj
uu8T5mCwM9TTgM2GKRJoArQ16suKoZu9Yf/3WUBobgmLQ7EiHRce7nRXyq1/42d9
7htVyAMJVOK8iV87YJsx13wcfvyxM8LZp3O35gre9tkSkU13JEopdqX0UDa7mEZl
Z6OJEra1sWVb0pZBcDeTNJkJP3KhCdLOjp63BGCM28EspqxW+xUAtXLJhFoSPJLd
vKhILT2dNWsbw69zux8bMMpzH9Gn6Z+oVLa+ThNrOvvq1IN1ZZ2qPoytH8Zs8tUi
994otJIg8uu3biTh1ou1HzTOdBzxZPz37sow91Rb6InMFOh8mnMHqVUvfWSFJ9Gq
+wu9Y2rHHq5Q4aoltgkPoCBlPcoJdNvtviU6ipp5fkfuaAfpmbgJzACnNrz8PXrw
RUaOWF1ZNBhjszPwMzRR+0LTlGmP6z+JB8w1CybBjf1ofclc5HKt1YnKRWXBRI/8
M9POwwvbGqX9sMqxHqxxkV4NWvYHVcGLrHYp50X6QcBd35vuZWgLOec1ruUOddAz
YIszXIfG6i47gYbO+0npUtS4ReAohnlHxxNfbsjzU9l/KK7vBUsb613eu8WAwZGd
c94o0LcPcwmGRs14qYzE0K7NJbjd2K2lrYIIm/byaRe3CEz+iM8QCxumQu3jItUe
Z2+xKyl/mdo5AtfhpWpvzuoJVapLLXW9N/osyJEDOMEyabvAV2g7Gv9YE+WbdxPq
PxNHnIPyvO3uh155NuaKRbq58XqNi/5VPQ4XajFNFwwZQM6V7sddOvJldN1kUqRY
jpJplkrnZ9YPcCqavTyvBP2cSs9pI9WEYqH6ZFpxRxvriwjTzfbNzecZ3zd4MUnc
j2X6Vao1JInfbiF53uIWWiDmmPqjo9A0bzkaAbk+ZlQ8KUg4Xhf08EsjZHIaTPAa
BOv++eh41+xWSB9uurIzjMP6fnMuw3BshG+zFbpNmRYtLmS0n0xVur97a2z1tBk1
PKbt4akNeFLE5Q+xwXow6dyO/UU3yHpa79QXMJ/e1kqkSdvuyQOZlvQIjkZu5rr4
q5RonkZPspXFGepSr5YEn/yTnTVl5zQnBCslnPA6Tu+OHgZkYWO5lf3/H/Tu+net
Sxv2I7GJrAVKChr9Fn9dOczRYcRIz+IL3rrojMwG49H3gx6IgIYmPtqlguJ8AzML
ylni0h/H0XGnHevkoepTl28s5vf1yuzU8BncBeVHTpJlr/pgVdT34HGWUQWe967z
yD2PBa16lQfiJNv8diIwPaYhB0MGnk7MdYHy+G+de+VkgmiuERHpxYwkWycO6UVE
mUZKTVOaRopiBV04aVs1ydsOtTNYY4LIh8Kk8sVQKl5RHvJz0BdsAO8vslol+5ax
xkvd+DXJZy5dpxdNC3rCT8Hc1rAXAhbqkM5BXYntZw+G672zNnlszFPDsTGlKcpx
YLdp3SVlPdtbJc9+wkkLZBQydLWlrQX80JpWiP11ep0D1t37gD5M0aX1hOJRK7dt
1B+ElAza3OUApjflZte9OtRrugzNLXa4Rj11o9E45U2AhyRo5Pm56ewtFqHkxZzW
DZtjooSPOPibSBAXZSz0WnYH7pqJXuzruWPgugg0VxFL0TwOqz3njs2xIPiJs0A+
VRLhlBoaqAzZ5mZsmeP9+xT2stzkGe0xK30T116fRckcxdhdz9H2gwgkFewTJ6/j
wZqdKvK1dZCkHOOImWmRZwf1VWJHV6kRCKhDcD31flHEE0M4f0rBVOfu+p3yjrKw
suMr4PEkbpQ9XMgV62Ac0wNNTHpYD5zJTm8F3GipoLidCykG6T2cgIIwBYXQHzQ7
qxMvB/ni942p9XWpIfSAjMW8kS6FRbq4y27ujieQLKlO7rDtGSRe09aWBsKT+5QK
aRYzRQ+J21dGk/9gWT5OP+U9XJV+Nac0dQ0eZw6t41hAqQTXCvhMTC+eMcxGGeGw
k7x/a9A4NeqMGGHEDKatqi34CGX/v+SqafQPBQLGlRIL1RUcSzPjpt8ngs188exj
/ulxwnxrtx8/ANtYF0FroEhUIEKy8+YKhjGTOWnIFjAL5F87sjenaKEE6tyLS0/v
vNdcuyqFxwhqVM0oWesqR4OiDBQPTxruYyKODMdNV2BOMjJeFdzvjI0xbGWI2TMI
sr/lqHO4l5F0VSgwjTNWY+y5c25Q0VMrgscG870kTly/UtcH8bRKhWR7ZH7qYuQR
EI9i18MMe143m5Q9YuQW0KP0Og0LGoIA2xFDQCLzGZilhb0+hQVKATLzAHSXoQ3S
AgbIEy94dhPxeagopwgm11vQTcmj1582Ljc5oNjAnNZClAWov5X8vJC7eYM8/SEm
1G+mmyKdVkYm9QUG7DGQ4007+spUFiheP4+L7c/WUs5kl2dRrHpcGcT/8/nA8IWu
29QSlT2C5MGPvFGLw4LwNFcBCkogh/2n/jA5tRFyLD11R7oIYD4WjaI+L/zm+kvU
1A/gLqZfwj1rjHLibyGzZR5yLmZj/gT1ibgXqqjHOkP16m7i6IJ3OiCO1KirOLcB
5JX2GPCXYM88wn2dXsR8cC/utGu2MAhbanH1lM2rA/TMcRpbmQEsYNNJcoBZktX2
67oc48fyBs0+gHpk9XfiaGPKmC0VRRV1Zhe3SS+Dw2qM7PlO868IEVY+XKSAGisb
+QOwfKQzaa9OboS7xzNFPXTal4itNhBE0bH08/9ykJEddA8ofS7yRKROwXaWc/k3
A4dx95BevPX+EpidkrbyFSbuyUQd+YfUweAGMA1dpcF4y+p1McPy6ChTqcLhw9yZ
2AKuwse9kcnRs+w94K6r+vmSEhhsocNDr1Gr/M6ATMHosNaI3S8mwShnplMDmwTt
I/HcajdPCUay1M1YqLjq8mC6lU790o1+H7zthpfQZUlrJA4tfpSa6Tc8RnZYdgbW
+XOW1UUqqAzz6kaugMp52BlzSOqKwiAvW46OqYCCTOkQHI9pFZ/hm3CytBoAdJnM
qKwJR8IVJ+6mYaAbffv3wxTedbXUaG07N1EoolSZ/8hnmVIgXx0dIXBF4ZFCFC9A
QxKVS9mqmKo5k/8/ccHJT1IdlU01Zmc1FHPlvDyZvZhNrZOnOUII/4DCuJg9epaK
lORY+YBcumVtRv6wU9ZBUD0bPF1TAaYj971BnbnBYClNH5eUdTu0zoiYuexWfWTJ
G6Na8/S+aspAxmZFsWZFY885NITSjKNYDD5BTooUJ4XJaJvTCGjM2UGblx8B6dpO
h1kf98fx+ziHHCVXwiVCgIhsLutzf2PKHvNAhKWiyDtId+mXOhSgL/taOysBG9E5
3DXsVcjrViNpFNKVXdtZwZfPA71JygM3zfMzYUSzWizLs04v8QvUVK4uQJD3ObBT
JSV7baXeeeClpmNWUeMtVN/095LdU0dpSJ+/AOLgKU+Hz4bUo5loClDJKdQilFML
fw77Srr/YxxfUKpekfPeLj8Tc6ONaH8eBPDdP4SIQPnqN+CPubP9SfQv9Cesq+JI
mYs/EC1hlC0hk4v/BtfvwvPCeG4VHrThV+ZOH6S52EBv3FxRafWhUfiP1vuiSbpE
ZWi+XNISIISUzibZpzmeqmArtYgxN9QQDA5e03nhPboriuk72KbqsKNwxtRDblZd
wt0q+vS+b2le96uHQXkCtxJUvNwvzhilkYkod/PDUCsmn/OIQCQrgjwKgQx8Juz/
fH15wZnxRzjOTy+46fm5blNsQy/R69t1BHxL1mIIGG83INZUIHCuNnkVSxYWPHs3
MOCTSadjUO2Vlzs+wZ5rkLELMFA9HdNNNWhT2e6GH1tQuxxkn+yRGt9dLE7evbqH
+GIoP2hfGimemDTv8HImR8If5uwFmKcgS3R1FUI7cZN5gd1Q7/609oVhwqpG5AOP
ljranMKpMeIOCmczAoxM54DS1Cfpz1C1yzBrENyDfJingY3ooWuc8WFJcrrL+D8T
3A3XJJF8RwC6vDREgcxTSqUJ/sxYYo/jxLUiW456Oze5gN86wNG41+ojvXigqTEY
T1pcrUccNbEt8NrsX9y3a0VTFVzw2XMQTw6sQrECfYmV8WNmvwjNddp/v0LiPQ/w
/i1Kw0NP7A5lkdA6LPumlEkoLVHH2PPd6DVp4t6X/TPSHkJt3GksRPu1ncfPovoy
5sKiDE5ZsK7k0qrTGhLAvIc2P2MxGInv+ds54D8gwZHkPALgDCTJGa7vzpDTYqZ5
XlvXQERhPOSyKH9aypEnfkVil+NR4nVSHz/+GXLmw/o8Jeghv9jfDgzz+/SFQksf
6estQ9mohF2KANQxw36qgW4d9SpB5TBgzv5dFIIj6EtSt1MHxsjb4B/F8tbxYpKn
AqmS4+KxDqbc2iH4tCpPWndbK1KBPqWikZ5NKekSb6GFG+TB4In8P5/rhjBase2v
M6k4ndGIGVSA1MrlQ5wUkffkZ3VFMK7U6igx6OlYIMHlpL/aHqaD71E1ZagTT6wh
Pmcd8/5CLuV4G0yYz3RHDP3dbsHfz5S77Yr6pmCWzXkBWwowSBjRQP0f2yJFmNLo
tC7vLMT1Kr1Bth0BWEU5KauEBxhlqbxCwtHObGBnPFFYsfA/MbAiKIzcqNnh6f+A
sqOXyNXv/4l5L/xXPzOjawtpgnB8ZMdZ708e4MUjq3/Jy38iPHV5k6HZLbuFf3na
2WWf94nCAxR6v2UxHFssQsaEEo/Xi2fUWrvd0svnC/SiEdwd8WE77nZNdJFi9Mzg
tEG8z4OsWKg82hyi8btkQVafH3cvZUA6YmZnXb++sJIBpOjGoX3A75fmapVwaC2k
6erUdLti7gG6APA8wbVfMyhly+Ldczsnd2tT9/yrjf55JlVcg0kBgOlFQ30+C+Nj
NZW1NcgTKhm/hjI5myKs1q/4hVuQcM3NzP5g9v+uv4PkS7B0m7z58WmwjAh5K8J9
WMb13ETNAZ3//F045pPa4iSz1d69M4bEXYbeEEyaSZjG/FKPsloe50xspHm7hiTr
9fDeemWFeAfuW8lAQLGsu6iolu5WvOnTHZArraOeIxSCUdViS9ebQtbiFWaEEp48
bH+WYecRdqXDu3BxHnkc8/ULFpIrfyyGL0kasGHN4qvcvDWIWp+2iYcHVf5Grslp
Xt8IJBJiedQcrXtGCb3iJCBoNiKoA4cgzyGPza/Ag0qJPatwZ4hsy93PKafqtJ1A
EK5U07FzOSGRCohRYySTk7r7JP/5o473zQid1SBd5MewqDuR7hCqIFOA75U3laAw
jdpQCJmwFwjOtQ0LLCzZeXJYof8HMP4Brj403ol/UdFZASvL6sNSEhKYyijJ1qtW
xUiHR1xGDje9hIQkvVDVLPKovna+z3ujFxXCmuIGiJng3GXz3bz2WERcHfk5r3rN
k3RcurI3UBaaicAyKiOtj/W+HwnawNtliC0CzDQfxlBzyVWADeXsLMUYeRt0pau+
kHeLawzxVHKauTKLbxgtxb9kSfj3ASPApUvp3dh0RaE3+QAW9qej5qX4o4sYw5MF
vvDYlQ03uAWXgOR+C87yc0e2kbubgM/F3pzqk01mdceL8c+z0F5YQ+Epq/uT6FOi
L4Rnbqor2egDMu6VXJAd4dVPTVDaX+2lUZQluxslZo5alV0Icpzu+9MHwdRF3iCq
eRU1gZ78ZeTa8uLmXEbgeQLUAjkt9/Vhueqyn5aprgf7saefosbcU3RjjXzBiOT2
v29su6nqWOBX/49IKz0mNUPAnNaC3xGxeQ/8E9hlUs+6ET0rBfLr/L+9SQW77LnO
xlRl7R8yg+ShIlN+Yds0XKA3ePA8k+Az1UX1/Xumwt5W5pqkpmV5YN4bleiKScF3
noMKtOGsUyPgMi0BWJApvFP2JYAUIoynTZAxb7sgU39in5/YzmKeTqBwpvikGkGs
OqIZ03FP9502WuXT3fwsvkJy3K+Lt1absLwF8/G23R59U6jGwphKwst/im+oMrlU
Iv6rNd+U22KtKs/Azlb33TAxSNWToRgOcx/2dXcaZugIOp4enuGusR5+ls8HktPf
/R/8lzqo81JN6NzJVqFgQQuv7Oo8GJa0poiI/m0eS0JW3foE1gZCxYxmDRikRL55
oY+s0i22XF9EGGA7Wm2C5SqcHfOW0dd38PvmwWm5PriuK6q2ziiUbpukuR3f2nu/
29QWuHaxBbpwiuCYrrDC6WZlMb1BnaWOLH+XN1yOoS/jOrbHqIe/lqZRTGDi5Drb
8p3rCimaoFstD86N1EszpyZmeVgzcTls/yK7cdJtaDHUfglQW7B+M6LrUz7ss+rQ
EdOF8vV6ynlnNuKO/arqAY9ulnhkmvyakG/BUJYo/o6lwVVw3UaT1rLRHxS8JHF2
5XLXILWoruADtpq3IgCdBfvEd8+Rt7td52ruoia3QY0gpEjG5OEtcyzHGeU/o7+K
JncgCN9InhI8l6ycPVkIwlEyxvG8qVSHrkAvh2GtUpZ4wav9x931d8d1X+VbhWD/
bsuj4Rb9gHJLZEe2Q112jAYoQjRDyTSuXwbunXQWUVildcCO04PE7V0zuu2/Boqh
gdIXsjkBLeD+CrFr9v3mqrjZa1rGwdjAh3FUm/Peq89VXJcAGM+YI6u14eJpZctb
Ze63Q81fTdPTIEQ96tUIMMTknHGOGsHX4S8sBXU7DlhTQRl2b1H5Pe70OWoU5++z
tz/keVQPanQxTXKVaKKzSFDa5OxKrNhGOnqmMFm6UFtKvK/iptXwiCIp38jxnxY2
wzKzxaupAg/xdnMKzw6BKXAtQ+bWYQahMVRUwMUQIl5cX8Bil5WOWuojzdSumqc4
+jALiAuEirWFx6pzQDjE6pBV8jWaTEV7LsHUPxMk+W9Wunz2lB1jvLeaERoGOQeB
1cRYLL3N1l/YuNxchujvUZ/UIgp6NgAFrPdD7+wt5xBecNGl8Zp4uHftrxbAplP/
6aju+WHmcWlxuQf1Ch/dp+WGUaVnfw8JsWt+XaTtDRSsOMvswCjMy/Qi4oa9qHfr
+9MZzD5Pr6BboUMEPsN2Yrm3lXO5YDdPspBEXDXwLmLIrkVSYw59FjAAzKHGEBva
8zMQJUOtadDafkRbkctfJTPB0Ag1TIODte6WO94Fwmoo59Lu8IaXbJKsmB4O10Gb
k/FBxlQS6P8SqurxsEknmEvHUdEBwgDhxx3bfgsOxdzVpR+bCXil47W+bPynkkGF
hS8FNDH59V2i81Pl9ZPgzsoEJ2864XFu8gBfH1hxEexOukrJNY9/IMv1gZz94L9j
FmMmUqQ4a/yPz+wXFG4OAqDkVBBXBRB2irETw3GCNGDjh8+6qwKE3gsw+iv+d9vp
1qv2ilHU1/xITFDu+YKCtr1HvGINshjrJpoXG4b+0XQl9CeTC1893LoVEM/bDESd
T7iBxj9asUHpQ5tvVxBV9cOuw4iwB/NXMUDtm6FtRf/lWe0xlykGswAGiz6424X0
qshQhet9bwYWS4WgQnnd0A0lRgFpcWL+HPoDnvFfBvOHRrLGSyVlhX1N6omoeEiD
ochmji/BxMZN++GYwP0tOqbfr7UoJfRUm7DThyAH1uLz/glv207R2VK799lQR/S3
Mn7BIjSLNET9il9Q4AdOIa8BRlIqnlxOojDJA87CpGtceSOB1qt+MRvxxk2fGUhn
Rm+p/ScMT65JgdY+Iaamho+BJG2jaF0yBPppJGNXv898ARTAvjZ01y3EBHXo50aI
hWsTaNxZFhALKOxUhVVr6cn2Jqcf10RJcnWXpJnsDLwf9ycuvMLmafQvwW5ioMlB
Cnge0QY7mn7L1KoWHmLj03lfLjFHJlqmmjZTGWL0Qyh9Lg63d1ehZJM/8mIjjthP
5sps83jKfeRxSJH08qlpwKNddHaVPKHgU/koysDRLN+byByPtJo9j7b0TvkpVK3O
fcB0MyvvNdIrKlJjHRBOe2veVQVgd2LuAeNhVhBzRszMQ1RYXO+UfN5LCPsSQ4P+
DMAM2Lmwfg4tSntBzabyb0EUI0+OYNTL/GuT8f2b4yZ1sRjM0pGI98oxFaUGLWGA
js9WhkXhR20rbR8gnLGqBnMLVuOzsKZqisvKF4Dsk3oL92DAg0Zug/Inz53TF6zA
F/j0MEtnflagKZ0EnmTSQCr+ElpNkogFGqYOBEpSy55Ev9MVbP4sRyf2rHppXpvj
n8fiQZqHUD+EPjNIiDJU6QvWHtrI/wXLf63uZWSnO4Z2K1EZG6x1MGZda1NgwbxY
kq6VxK5HaQ/TBfGfl/MNWv9CEI7R3xxqmgnQokKfpXEzc17gk2AE9KV5VLCHAUks
Gyd3OxeQqCCkmTjOBYTxmIjkb7UHIcxYdnmwm+AA/aJHgawPbivDwCP9FhUQaDDm
/TJFxVd2XdaDoiM5w/JgRIGG27xBmO2ZO7BQWbKSQXt7i1V8fpr7yLQ9f+U/T4cK
X2aZvCdwkvn925UHMTnqzu1PgBCMHbb9S5kjLxDDhPR1fH8WnZA097uzSjmqABve
RtHHZc8zCsmHh11rvUTIb8reWgZ9zEH52V3r5UuqFDLb0ZpeZhqY/if8C9KbHjPw
88O9v93RwKJcDJbiQLG58KZS0H8t8GQfbBlqWw4Izm5RnnABAHNKiFd8jUviNunU
SgQ0cnVepvX0oObHFRwcrwWhg8enX+nj5vbWVQGcskGCfzYuZChogR3EovFfUnv8
IV9hFPTD2klDeBC7DbtbkGTSkDqc7nxC6rtH2zyGDjj5NvSivNPh1uQp5KMBI4Dt
LNMJopbLEsG2FabPAOKCkfnK4mICGE4kQXi2LQKQ51aD+HDNSEvHZ+YOeDFEsRIG
3l+hQtn4ik5euc3CrJ4zF5ZCk65TCXnws8ZxFvQQ21PFmV2C+7yHOKYKBDa3uh5e
Gaa3ykn3lj9S2zD11ieIUN4Zyr1OFn4dluxVDWHRyghD6nHfZL1NkNx5psWdNjfv
UK6AYqOAuRRits4YknaOsdEbnfTeLE94EXFgb6F6i3m+Qu/PvQJvqaYNWGn5zECc
5xUQN69U9LFNPBheJ0RGmI/XkbgIgbUPM0nwUD4+ZC3BToxiI0XOLcR5n1Yfz6ZL
1vbWYQlwy+F7TydZVZpZTueI+m4grP8b6t/eGa49jorVB16d5cjQVbARhJjudZ2H
4IfwOGNIhU+oqpBqQgjcOXhnq7nL5t61iK0oNBD/vqrO7BAptaZkdjmWiLkcYNfJ
DYXJ9+av0HKIoB2o/tV5ddqe2hkZFQ2F5Hdd1BxndD5m4Z5h2g4PFruDPp8vvHkr
6F5C0MIX0gsG8eOLwVAJiJAMQ3efZyv9Z7FoYa/+6KuQ7DSmklzSq81I3vvfdpno
R+Y+wzNcupvzLn+oo82ImRynYXcMreTyb1reBtnN2/AuEZLaYNysHDB0GUN3I0Ly
C7LwX9AZXdCEjeOO16rBn2SgVCnCrVRCUvu+We8Z7G1sm956My/BagaRZxMYTBZJ
Wo5DJFsQyP6HaBmeVkWyCRjJkxcVuH+JrBCMgXvRHYPDvjosBS/yNJiFT/0LC1Ik
evbwrBZ+VsYsgb14h27pMLQn8OvtLe0/XgH1YeWx21XltRlyMFZUgEt9CxQwSKno
YFhe9qPE+U/Vca0DoQOasnsPyACkCi+KexXycmWbIxtHnN+AEAn8zx1Qb2C10il3
Q2Wn4Ar7qPTpB+gF8LHAWHacBZa+sW3qUMLx0cpLyAv2OcZYEldXEXp7fDgwOaeN
iftLcTTfHIigkgrTryAKmUOlmzdGprwfNR25GWrCtmdXl5ti+4bXEC8XD3TX+9DN
SRGACHZTPdwxZ5c9NDXyBxrSJD5zepIqsmdqhP8hNwPBev/Q2RvZIt+kTcnt1tty
WKquIkyxXB+GVbJjE5sEE9VxdURp0AaXYcN4/kNwB5tgL0/8YDBTSGJIPBGGSk+D
CC3uIxsSkTv++ZVr/3UWPfaRdpKrR9PaUiPtuCMLemy94u80NGJyD4RGAf661bGg
IefMT/4ZUKxpIcJCiyc70+ekkDvuyfh4VWJRICnSSGuXH62Ayqa08LehhicIkUEG
h98ay0IruNWboek2kwQEHhUMIowwHGh/NxxtcOKGZBWVb0wewx0V6rGmMyG6/fzb
slt98iJ6Yqg64Ciwbncu0KE/dZbLd641Vk8DyngUrevpUe5soDQlij8PHKZn6Eub
/8KntVMciTnrdEYQmKhGmG3Ua1mdZSTxI7aIU5cg8uWtihhpjfB6wNOUMTnqi+mO
bJn+3mV6LxAt+lwFLiHPtwmnP+mwNA2Qqb7ZHbSAf2wdI56sGkSk1mFeFLps/rMs
YjOdCqYxZBVl/62utHR4IMfVEOPhNCeSczlbG7bnmgublFHP/SQ4gojVVBa+ALSj
1GTTJ39laAJWQmFD8AxePfoqvG60mtvekeoPn4IgywLAWkeOQ3+JU8qoDjBbwbio
wriuQa66C2q9LW8GOqi66xf9dZgoCZ57dSPpbjBWKsMNXYL7oM0DyeoXvHxXHS+e
ImaW6/TSAxRbf6t+iDeY8F44x+B47RxvBmQzsCJ1opqImDsEoY2ef+6xUhQ5qO+a
UqUnUEhfxmRT5Q3TzlQZMrd1f7V0TkLEvrYVreuTrEqz53Qhdt7fr7jSycNzmQXD
uMYsq2aeyjObtF2Ly2CukgUUaDHFw2Q0G6XCPSZZ3PnSJxb1tpkA8x5Q/Zhj8svb
sY4gnMbJ0rBbtFq88STYKU6UEM/LFMceAAZNKPEko0VR3Pmj4A2CZ9pq3C5qkWMr
xRFoFbjmbwLwnXVj7NQ4l70h7z4QDUF7npmdSVx3j375ImCAuVovdjTL47qmX/DO
t9P9uy/A1bhfB1fnx9pzQpGloQVfiSvb5dzL70RgbTGaOG4P5FpSlUlO3RjKHXNF
BAzB55t7D048SYuc765LmSRsUZsk+wEh8nMW8ett3HSlYxOe50nWFy5DdgcV31Wn
aVTAfqmUujAZ0PWjcHTuu6wUgdYS5KwLAXQLDwiZtnCje9K3/pqj4QgFvknpgB3m
Rb976pax3SuXu37VnEb8FO3MoSlMib7UjELosYU0IjR5G4vKnKWHhd9h7onGEdc8
k6cYonSSmOSvSIEj4ypTsdVND0Ty6kOGFHWxKgxRE65/qH9dHVtyY1IJpMU/ZN9f
aK3gH3LDdiWiV8LI8+ph37MFH/VulV2R3/u7YeOgYJV5kACGYM5pl6NtmiPVg0RM
3hB5HtF8dfxlp/weMcFPYhtM/xP5qMo8RUwThCqnJhdlMA+99dGSVT+HJ3ri4M/k
gZGwtTy5MgoZ8fVAwGi60XHucvXgZgvqP+vKCwXT3jalntcN2jo2N0y2KqwSklXg
KCSi5W7bTy29onKMHAltP1er/Bq3t6UeCXkIDC15joWaj//16gdgofgwn3N7JwL1
yUZPXM8d0EQV2iU7egnzYx3Mttb2WE8iEcUeO1p4MDfM+Vlkb34OLI5reksBDWx1
PpD0ZeXwNkc15Q4R3QeY65DT1EdAYiNX2AhGejKEZfNxPeVyTaojIHkyGY41C9ek
pNLrBg8GrNdqdbOwfZM/rfIBfjbJyVasqUhfXooQywR4xVLd6p7YQISpu7L4c1uv
+1FpSDzOxBdb0b30RaoO4Uv1mfFFQ+TWyTO0yHESfkfkNhWT+bBSkm13s+2Q0YM5
OaLLjbkKkqjbWXcWzLQKogpZMuXLB2lVYHuEwsbH7pXMN4ooNr0HagM+QhOLOSpG
8QoBdQmB2NqXnvg5JrFCHm+XzTseZvrDlfmsH7GhZeOYdHZfCsiNtmGWQ8QYO/fI
FdLiY3rWuWpHA9Z8t3GrYN6KK6ho7GrzediAuz1jSlOtmAnRQfIrIgVlNVDH/KHD
B1j7BJJhKrr0JtdzvCOkfZkygT17r6CFTw/+nnLoynt6VhsWe6CnglHaNvDxypIs
CeOIkjAsc97L7E3OXMTKZwk78w9LaUoxe72vVz98mYN2FSJxHAuTpovKhphgcfoW
DZ9Ne+VDT+g4JixFrD27StONIGCxhA6LJkbgCm31JneLHU2a3EqdSuONAcWyrC93
3q2+3KwhwPbC2oZxSKNfxWQnccyS4ARi6LiFZnrqnNu76VdvhPPnpFpvdcMq96lF
h149f1y3q/jD2//Zb6KqSv9xjWFHynIieoG4AgxW7j/nEqxYyw94xS8BFPfVadTV
f+OBdLFhHoYsMXAM/GAnxBun1p5FCpCSwm3u/d+cO9GY4gZOype7TVEhff9WYcKb
auA8YP6czCPz+eW61P3XWoyjVKGSLJudrN5+RBV0TW9U3GVAyjdwvRpe4pOEszfN
ahwwI42mu3r9POTxktim+0H2kaKC50LfCbxX0ebptXCjc2rrUitZxTcbOYDcTAM8
RdbE6G+TreSynf8loz+9O0kxGzlbvGRlj2xojp2kHQandTyZNTPwYWQylO8GXuLc
Zh1znyibShwLcsmTalRQ9tDgAOCfH2nTCGjehYfFTpkhBfRHYpjhx1JDjUqOYKTI
6QxJ3f5BrZ6q4EPlYESDP3RqKX6NOEL+AMWlAr75xb8Wnin+R3Y4sdNCUq8jgpY3
aYYNse/KLOBVqiiEt+GBZ7i5xPHP/lnxHDGkcL4yMsDGu4r0f72cwg+5Ooy9qA8j
THwSBoQ0hRBOn7NL62ti6p61PHP/kSIHXx37ukt0kyghA10YbFb9YYJHUiz3YjSW
b7mmWTvc86kC/WZX3nas+GLM/Ko7PuHYYGeoyW/JgWLNghTZrINGJWa3aEkwJWM1
RuJNXZVabrpx5uDwIcYEZeb2YCqZOOgC6O/LisBxS2/RjOB6h1YKizC0pVBS799H
Zgsz1dqkMF/alDqM84G5SCWubU4KVknbT0nSsAXgQHJoXIeP7e3nM1L+5kVSp4lr
xW5QLDj2HloSbR33Mgg+S/G60r5hbhLZZ9ggYMUahSeYGYPMVEj+/jcq8thY8lqg
4HYkRZg5CHrq6orz9bhh4+liV5JdqVH4OMdAKIaKHTieEwN2f4y2e3FZXmw2Z32N
dcCLPpmALCVBdBOfNnNN1buzFO0gB8EY3MFcNX1slYF49vCLn0BBZD0R7lwXbXq8
jgHhgAPbxoJzwBOsNXLz68OHY9b3cRdRXVKaxTIIpQkOAWTTzxxXIKXQoNqgp5u4
j4EGwcv6mU1tQNvls2z9qG4jU42UfJK4cxSC6Oc5FwdyZVhibVYPicOpOH9B+Sie
N2wTYVBjurEQOSqsJ3ChYK/LwHaubnLl35rms0jzi10bOYdjkYORXpt+RlD87Hwh
VNiUGBG9WK2/RBhj1vZmOnRUgSnBe2USK60+wLYsTgQ3CXIGGVsQTuxhfgIT4XWG
atCzpnh229P8jhTHTx04tKYKfWhbGNUP9g/hwzobZIHOtwgF5szP8SxZ97E5RqE5
ZC/rYdWKUPCGQWQqo1Ag6xz5ZRhmxtYf8E0+7iybEpTvlO1czMTt8/nCjt5rmeKr
+uRUnMl0p3LYfJcBCCeLDuHLQduR2kiI2vnvVcMs+59r0bszjWc1aKG77Qbqm86y
pw8nc8uxlDpeAo+rLIwFWFwHGjLQrFGwYq5AZJbo61dL7t+4plouasN14p4/RyvF
DLvWWy0lY5+DWJiNNFZwbU/e3qlSZO4/RXQvs4s07vHVzYDso7cbkP04rCB6mNCq
0BiD+W5+u1M5XGx89oSMh7ZrzNGvGqQ5czOHZ9xs6W/o/5Cz1/evV1gUhLNOSR4D
2Q6oLMfHtz2lpMop3/6JiA5KKorfIvC/CBdIrEs502C0H7dmRPHi/btaLm7YFcX5
zB4F/m4TrzeBlmbpnHfc5nQvfdjksd2cIZGBkySS6Z5zca8dN3+yFGqT0pEAfvpE
eymHGdKErnnQGwHbqeOK6MKSeKTxAt77x3NilaeHslY83TuXkN8pgUnoGcCaCy0n
yHEatLciWv5stDvPjnjLCDq/GYWOlkx5ri2Opap4vyjpzJb1fphZZ0p1zBU+sf3u
zv1Ow3Ft+u/LW8iI71UniX00SnVEf2249aHHwgg4mrnE6zHmgigYzaZW4jku4w8I
/jg1ZJqFwhA8nO6b9UVHaOvJzBKN/bYMTnMM7ZqGA8xE8K/Rv9nQjLILXR9fac0s
7gpQYAd8YNs74ghKLHCVv0+/tSb2fMQn/ZKDHFYQmla3RhRfZiELrTEF1qawAuyR
qB+lKmveDR5ng/rKiANjiBJmjwoGH0oQq3tQs5cl9iKY5iqGzQYTWP3xwfQQgl/3
afECigJzgWIKJyBvhv2SCP4zcposdnx/siIf3oohpmTLs1a1Uy/EOuEeOmgWTorC
1mfG9mLqTPs6ATmzlt8S5bOXZVSoVaJeHIeQKbZIEEbbW1SZpn5nWiOQqh2k40Gl
tfG0fPVsyHLSwTjV/lAhXYgh7nodM/5UH+r6Uk3Com/kjBOsDiJAQnwH8X9C+RuX
vrK5/6dmLWfoXLrmSsfQIF90yEzeTr3dQaRJ9m57u1zJGFoNshZ105Z65a8cQPaV
I2LEWgFuqPjk/gz4K+kh+80LgZy4G3RZOyatZ55pityLwtFqrOj+SrNVBeQHLQ9u
t0ipeMGBFdQNkgGYT5kfgB371unPr/rlPI3CMgG4pPV1ekdPS4A9B7A4y/5r2Y+s
hV05CyiY9HbuYrlI3ittiKOKZpoxFlFx9ADRLUqd9Axffx7ZleqYYMgGyP5EEc9T
7Zu9x+inZc0j9NP2f1FcciVQui24OlLOKXLtJzGkqJjBjhaD1W8lMtu2+PYsX9a4
c7cqdA8l4yU8iBTWaZH+/fcT87GxawlsQM+tPETLZywmCDTUfZ782a5t4eg/xK5i
BqEz5U6LTvRETJWYXvUrEkxstcYJfHuZmxjlOU4Ch+JclyCvs9ZF4HjFqYIHc3sQ
4BUeuRTXAcnltaoK+sU4qCBTZm3EIQ4lGpYi1TWJZ4kaN07YRcElGweclDJ0LMTz
NygGCgUTjmZxjtonqsN8jkQAvzUNIHqgj/lDvlm524YQrabGU1PHEMUhfah3BsSW
eb7O6itDiv/5vfzSGhTuzdDZn7wumvZkMeepqPsnjJ+QsYpYjZGBYW0ctCum03ii
vL12CleHYojoIc7ACD3uhj5SMkkDbf6R1Ndh1MA1EsSUpy7RM2VsMM0NI6tOmaBT
wkg5yAq+mTiMkT/tfE/H17RnqPT8oBBDDrHQK3JDghOcsj5RE5qJu3RQNR7hhWFe
7MirewV7BfGHQCjMzyLdqIscamXF9jhq0InNSsAgNDJfKsNU+4fb6gHszn8qYFGA
yC76jjt6MD9ZOZ12A+W34QKLlSl50LBquAfxb9KYgxU5JgDDuGzYqXfRDVoLcMzg
p0lG/0LLZsx3U2meN8PVzn9MSR8qNynIeWRebbsgHUfv2PPcHcQH0kDDQVJEZxdk
ux4foE43PFkWkyjfZbyM+mcFKUweW1iVvYJCd+cXOQBZHQXrkIgAt9N1ckAiijxG
OqK+dKMfSpujWkKlVh8cmspcGFgGrol2Hl70yjgFtWLxst1x434tehDvaN3gPJ0D
GGkgkiQy+30GkrrWjPGc4uxHqcFWwrLsZGgmXO988nSPAze4kflkKrQ//DO5m+Ne
rtwN9NiCol4o+hbgDekFjuetu2EKRMoDZbzj2PlAzfCswyi7yC61/iyZhmYPSxr5
t+bmy14KtOr+WrPrb7flV4MCLhDtac7rFgFvk2njccTfNMBwYhHt+NbtW5R/0Uyu
Il3CC6RFqMwArQW4+pDaGci7s0UaWUXQZclcIm3xT/OIXQ7Mx42ye1R67EevPIvP
A/Kjr1rx3uso4WAqohStSlQYJ737P7FJXlfhLSdUsD1+EQ8xDjmM2jqHd79bzLtP
y9CfU0RUbL9XCIohuqcREDn/R/n8CJie8Vs28UOMbrQxfkfCyCGfhBepTQw/lll7
atpQfep+fvv6966HWwTNUm+z7fTBy+HqtKHLulpNt0tBH58sbVBZrd8HtBaAfmIu
T1KXLTDm30Nw3gRo1E+Bqm7nYjcnnNQ8voD6kNXZShVBJrfiDxF3m21hrEDJ2hIq
iWeykFONlNbWdd05uxeTJ3rJ3m22QAD5bABXs1j6hDYQd97lePxdtNdZ52ja63j6
+PvgEzIAr2CWMidKI+sFZzFTqLa5gY1oha7iOgoSdOvuEYTUOKNUgMKLPA+oKCDR
yV5MNzfPCklPWIlPiA+stxS71y5FDRz3XvtFGADm2PGxAIbJR3uucsPBZAn1ai+2
APMy3BVzCR3FmMFYbER18lFNqOyOyZHljW+fnVxb1ADyEMXdGiBcJX3qsuBq/qnC
+cGhHDBggONdojJEYKmGMWb1mVrh9TJlvgiwFNWF0zZGZtdZXa80zUh2GfwtMXqG
i1tLt8u+yGPTIEsmua0PUNCWmFkwW8qL75Wp8eCYcXuC7pjrXNWrY7G5Nyhnj6cW
HIvZfcAuPyko1UAbFU0O+cysN+eb4eS51gicH8swQTpwxa3GYK7Og0XI+AuDDDsy
lN3lqu2j0ZF8kq1x/j0EIzYCCUrr3hTtRHGghEhl7SeLB0otPsKQSQld6Cy7brZG
fFQMD11oxZFsK8QBkHvSWcUzPaxkbvPD4ncfNW2JmD8YSAq1RZtiXFTTV6yaP2Jh
fCwzySvCe0KYzX9jUSnhRa43z56uyYsuUXTqA2IRlKsrxjdZD0Z7ebjSj/PSt/4z
zrL6SRMb+4+EoXOiW1EQ0i6CkOhJlHExi3fTet7sanVCHo3uNcBOiiyHDMDSD5V0
ywHO33ThlwcaQnfwoh9Kx0gNjBxDN+BGsi5lQMO0C1gA3/KiJDHYukoTWWwStyP7
YY+tv/dG8GEoTWaPE0eDyOcBtEizSxGvCggEfXu2YBmWmAKZI0xkPcEUl651+Umf
E7uDzZPwwch7L/bW4wesJNvZjlA2Ay8rtawhyhXyxQbD3jGqRq7CcGyHOqf/1WvH
9Wz1+0EDi+XRtH9h+ByGftAE4UFUiuGXbYkonWDJagVr97iLsFiQolRH1bqOoA7q
KH5Z0/3I2gS40GiMpPrRHhMvRwHPtUrb5DrXqGLOfHEOv7iFWUjcz73NsL/1vOg1
XggRK7VdM+g3CvbqrnhCFG5kD/dYu/JlBlo/2aCkPCDEUNKwCSvXOp74n22TA0ND
xvw2Y/GPQnanpjsztB1p87YYi6S0/kD+A6Byj7vunZxQLOh9blLCVvFxD/QExG6T
ECcXdNpw7oBI5x5uBN3yoYf+HFXN4rBNFWB8EipJ8CLgEUCDET4D3nfIgEeIZZHx
P38J5rkEV+4fYKN6mebgJH9tvy0qyp9MePElZnBqmunDn++GVXG/68IMVdlg1DpW
i9ORYaStA09zDvYQPRiwTZr+xFx9f+mxY4zMmhWthJnmW2qBzy0FgtujABgfJ4TG
QZy0NLII/kv5udDomE88PdkWbDxPki23UK4pbtxLkZdTvgvhHMQxRFbZLVG7WPhK
Oxk2xr03GXB6X1ZFcDjftVRWM2yguXxUeROyCTnq+CZ9MHiJjGZJVaphxbAQoubA
LLazbmcQt2No7FbYUQE9/fnZeCyUbKpYPKmlmDPkd+V+wGIEHjGgFpl29g0wnpq7
gi5PIspbtLM4D5YWnhVJNtTTmZebez6yXiTW9hyFZPCh11PcY3p2CL2AMCdHM253
YLfb2ejSVzj/AImGvuASdKy0UEMFE0s7xGsBWU/Hs1cvfKZYTh0OvGffne08kntd
ocxRX09LX7vuTx6d3cjyE8UQUYvPQ42BM5ppBi9EQbg58lxOiTd9M0Mn14NL6IX2
voKkj3ohOuGc9ON97DodpnkG3CaAX12aALy6C6ki+k6TZtvmtjlKbH8h+Xzj9bPc
43so7fEAJJA38LDzQApQT30WgqIp5cN3lslyAX+YQ9cRORA8tTWtSkFi/wq64d0a
aBG28m/QFvEJUKgmB2Nn1DsX4sLaJkSnoebiT+5tvAFZdKJTNkOkR9loVz0uSm2H
G61UtD0SWoUSsnLOwrzeYdKJpGeEqUJTyLEDbCBTlKKNnpKlzJUe4ETfR5XM9xrs
zKLZQ1UDyrclceB1HT9b6bPbpKaiGoTKLS1NjI22teXVyhDh+Bd5TXQJ0IQjegMx
5uQaasXLAyiZiatYpcjKR7B0GZQ6TU/PmRAv3X3f2VuBGK0TKRARwi60dv7UMt6R
0xvaMVY8vcsnfBO+AGhkKW5FIlte53xpRnONb8uFAk53xUuApNa6+xGb620nxZf/
kKQDTFExV4w4gJP7i9/ybin5UduHOX/JXWNM3VWT3ghZ0KZHDSwYmgPwWVNJ3+mB
vZA0N+2W5O+rjwZV+mDsezpUsZX5OPad4W2IGW9NHChU5e1gjY5RcFrIB5IEDUTA
IUyntKGy23N6JqhLEPD6GF/gAXFTHaDU4y/vjo4j6Rp3d5Z/kf7pPC/recaGk5wY
bxr5gAjPfdk9PopZbEqB4sk85BwPDroi3xhTFP6MuWlnvIaVmvG7wwd1r4iJ4Clw
gREpbtQlrQWVtfCFYrimmq574/MbSfgeGwYVleEQHJx2n0qgxI2jWy72haZDZSle
ol1PxtZw4Bfy+dKTmP33LOwx1K4M3wP9aCPNAmcr67eUq/vARqRjgG2cNWbigO33
nQsMGzeqjn6cx8+ThgCfilP3xkgCdC9qpRLJgVlajq3rIu1/KYs4tQ1liEPtOtsx
XSgnT+KZvIbGL6+U7ga7s+8EJdB1b21LiF+/IzBuxoueEPf7NWg/SAgGKwTNspxM
rc7qtMr6FMcTGDuXWMWLhNVQMVeBxjCRPagKzfD9ROOMhSmFuof3KOkBdFD4W1Od
Fwy0iQ+896WBPrGlBQ61T8M7FYCedQnrnz/aV34Grc145/YfDMB5T1rveEztuOIG
/dD8izVGXPZSgglzj6rgJeVjGVEBivAbdFq4qW/O2na7TfFbuo3dkDBQLC4kJmrU
jZFmtQaSIjzkwfzsgcGvaEFyiV8K8BAHCnt2oF6vZDrWQ0J/QTVrndyjXLeR752C
+33T7QfkVNehyDgoQ+SQksc8GtGYs/FwlE8J7Okap1Qwb4svxl4+LCep91bdqKat
WL9Fqxwc4TJGh3inIZZW3Funoz9rrKma7ePgHE/VlYRC4NeL5sGlLCQeQ1aN8t31
0zABMOoeReqYV5f3tQ6J8JIRQ7TC4jOCzT/6nE9RxqL/2URfa8EYd7B+fVuzKfxn
SqD2m8E+oYplSUft4t/wJNSYjAwjglxZcasv5m7rxy7AydiZ+/9NvtE2PJBpnDTC
R0a58QBUm1jk4428feht6pX8/xUz+av11lw3BBrDnuDzvu3arsLBHsKROfMGSZ4J
u+D65zJXYVEWl6qDqJJgXY7BKVHRQq3V/SMUOPT6NRM7+sVIWn9/ldOrt57R1aIj
ftDOM8pTvpvRnl2pKCQQ8/hgDsCgNyWGnIct/iU+YEPT1CGTH+hltTPrl5DPdX6m
MuwcruNHd1nNFnzecq2fTpyduYzF26gJJMhAXdW1hAcK7NRaCpvqyjcklBUcaIts
SRwyfQKO5D8xGdhD/qVwy5dyTfAo2lFk1EJj/5jETXGsqKxuR+sh5bveu/afrOjX
zmAzKzKwg7kLvWc/IJ64ZsTZOHpQ4P+VrU1G729BKd/oPshHE7LZyQRMyWZGhjle
2EODyLERhyRxDk9V1y01VJ4oac0s8hvG5iUoSUrYG5Kn3d9I9SoE/KqFBKlOtuXl
A2TSZOLvaZVOjALDSXVPpoEzsj+SZwhB9Vkxi3hc/GfJfEeNrHx8fN4cpJdPY7aA
XQ1v2I4e7p6dvdq+jKPiiSgRH6R/BPBaaqx7At7Vz039oOvvFEwBZWWyWFLByaZ5
9RclSf3xJX15QhNbMiuMttZW1cFYcLDvrak3E4apSUwjArrgQ1fYFE/osDgziFVn
RBhMOHe7BmOFOARSCthpyMDzFYSRcDGC/poSmNhcycPEFc5PnOpMgVjBoYNvMGH/
mnuFVuhD4YTPihuI9khFBIj7wkQ/SkHcGLf0IbBpursrGsDRkukIjThgWR0vSzzk
WwNQAAtcwncxNJDKo5TXomkx5ywmI/vQ5uAvnltd4gTyaKZeUQrvb1cR8zKzFpc3
RmNZJFpG3kOn++batW4rmtFk2OmrY5buNcJc33fZblpwTAN0oGhjTHe7k7CmLTAa
any7kFmwaW/H+Z3Ll3jR9kiU6O6khu3qUo73ojr97diGP+FkYRb/KFWmBQtX+osu
cC4DNhVLLPv6/nKMTt3X4yrQMda9suXm/BEEl2ll5+p1paO6JZjuy27OnCtRIMQW
Gpz69pxE9aPBgWEzcuY0QUrtfaosGDerIkBzhhzTApMG6Jae/t8SjcUJOH2Oyyyk
x/C40RRkPqfXvopX+vD72ulcivql07yJynmtI/lQ6PrSEJO7XY2kF8ucWwGL4s4R
47U7mPvKoh40qQH48GSvXzR+A2mRJxRull7bxhmFhZk1BwvHnPi3tcHv/lIXYnYJ
MBLIx9u2AKEcXAnw3DESSFAXLTLqN87ZJQmjciKpkV1W5AXkuTfgR2kuwHtDshms
6FrVWDNJHdPAT7n5x2PsRmqO1LgLPQNsXWSUTtFBRKyl2em0/PM5scMfAU30y2V5
XJoMvSee6jsySe6UNznHPbCxuyBSzApIQNxlArLkrtvQ5BdRwxb0veXhQAsKh2Vg
snJfjl5v/QyUe/KrEuVginE5hyWInzyEO8tOTl+fa4NYPoimWPslyvDUbLqfmZ3+
OrbEo8P3OPhl6OOuU1WbySnPOPMzmxBZIl6EuTsicMYxHRWBZZBYe8gK9HsMBx2e
PmY0bLZ47kWNtKh7OPDhfAHYYhVwjXxLY2/4+X70GpDyvuv6tB+Zc5F/OO+2jS1/
m/mbaLFTLQyAUTAVoGgkBUunD+gtOYQHCR8yEG3fT7K58DZ5Xj891dwwB/1K5O14
DjMrgYh9Qse+8M5qkidq9yD58SmsGIHgNftExVzsmJDoVp99anByZf2DURYxhE5D
ohaJ85ROP8d0lALWFP9vtbbsFuHyopHnRQ9acIbVY1VmYdErpeQN1u1oZcZT7W0N
DH+k1e1OgEPMWha/mPboQEvEZVQzpSU4EvzH1ENExP5FWUXTAK9/7uLtNygNnwDB
dpfqIlY9NYKE9KjGmbzVe40Xjcir8h7oHs/DwH5bTjw/MQdQLL4bNGxk/RzZH+wv
r/1GK3+CCSBpfcQEeG0YpILdvR6ZjUU7fOqyXcSaMy4uA3mA4X3/1fH2woKTcQI8
MRCkd7hJ0tgnglaJnE+eJT16Q9Iachzj/MNPkOjSNSzkhsoQ3kCH28AU5rFIWQYu
jgTP5E+Ywr+tHuRlcc8/b5BytbA5ouO1TwxVwFwWY4duX43dbk+5YXI4FaMOxtZy
JCH3FXw3Fsg9rQQQc2VFVOjraRB8vtiTkOhEk4HHq4RKgYIkSBQraBuTNzbk8vO7
/nvD1p+1pKdnZjLMppXicJblIzi7APiVXCspbyEFJNpwdDQHWcA0769Cq2JzAsDZ
yWQMOblBOUpNaqh7KASw6wBoCbB1wfxNNSV2wBtggqY8lO+hWj6bHag/ZW29tOJa
S2WZ75qEHCK2HFuv/+ZrOfVUIs2ty7djJDUC4Z5bUtcZPOVvrSKTJt14VTugYDiz
BD3SCdNWJreHxT82tF8CaSRAKwYmuQNkzsb+kvhQWGjsRFVU8JjUK+2ipjCn+Emj
TJVdTWIhWHycuneZ8ApEyzZB1Knms5XJfNcsHi/huQtKVCpz0K0QVze3Xf+4ierF
ORRgqOu0TmVGLiPN2ZQcaOGN12hVAFMApNDLZPHK7xLeUwlRLkY3nRL6KEvMTaQg
goUCa+G7IvriZRCiHyfpRWuaYQF4pkJzIHDCwyITLarlDE/OZcH4UJoXPjGmCQZU
R/3X2LkIKvXlsNzEXD1bhOX79PmmX+5E7xjBTpN7rmG8fimw51qcHFbs4q8AVE4/
ZJhclS1XHidpWm4q275piAilDK2qaCPJ2zm0TDA+mts1sbLY8FoVaXARmj3CBJSs
FgczeEGRA1dIAXZNx3lprVxZgj+1WFqoHiJlKPDH9ejKfd+6neXcUQ0wz4QPWUl/
RplBZvEXfSP2WVlg8qMzhSOaN3kqUqkzbLC9m2TACFpLQAkpDw1VqgfBk1IwDsYY
LxzsmRUKKoaDWTlmZrjBWkumggvXid6tpOuP3gr3/ceuMMSZgY7Wm7h11KI13Hx0
hiDrRzUMQHdJIe7/PNtgYV1GCaNKKe1tVd1tnrGIO3AmwxaUzDFHxuSNsD3qZ5yu
2xTr0kQinf4G/w8TPO1dLkPXmABwrvhbT6YHlZ8wSdr1cgUBiMm7stVKvjWD3q7f
5mE3z6yrQIHkvpOIkYMOYSjIw53p6Z8XtBOuL55TfSv1CzemzzrtVPCCk8zbivtZ
iRN5TEgZDJadnseOyaL8kwbPKg8J2pTqRkJL/jlISZhAZpfdNC/PYLc9r40PfCqf
wc4vWrsnghTkhnvqqddKhhq6p/YKrDKODhqMu0ethnnqyZ580qan0LnQjsWK1OE2
WB2hLnxfW4rFuruPHFdMZmnn1Ust+Epa0QC05UVmxAVj7bR8f2S4Y3LB5JogxkRF
TEvYYN1NAEZtN5/aQTOwJxcDrh1jtsZF2GJ4HRqd4likHwsQFwtEVtV8hQ8i/4+J
tFrbROT2W6nCJcUZohhROXzapMSL+uMNXS3K/Fq4SV62qgWewLgKWKtZv8kNhb3K
wd2WliMhtVNINrrw0A7dZtHgY+k/0Kb8feDLayrDPz+vMQ7ifHeLhp18FwdaIyzD
Og+1PHPqHrnzujZjBPmQ6KuBVYAst/lrlLiRhgrHKGZgiRyRPGajny1BZxg2vwmO
xTgwaahfwz7LxjZyVohBgWn3zxPXmKddqRI1huJbUDQeF6KFQXBHM+ePOntyjIe4
nWZ3JEW/W8lGsUfv0btzY/JwkZ5gQM1sI5fwWk4IU0uqrm94sO1T5ItEIezXjfNI
ORFntEkXVQZKbyrqbR2Jv7WiRlrDqXVzKBH14bvC5QCrOC/dWO8/1kojaON6RNIi
B6mdW8HvOy34bYr43HLaWJZ3Rlt1hoD7LZN1xGR/fdhc/gQtQN9bEpOTIcsqGEyk
mx1Khj84WjLGICcWOpD2aBxNnshuIFwS/8XaDtaky4T/d7/8p3n4jHfJ4HBHza+V
alzmEJFUQyCn3nH/78RcLTtk7wKSHq5l6pylL4O71V0sWd4nnVQXsPd6HyCdyuTA
lnu3Cp248m+gE0QFYCWkSmwaMNgFl/pCuLXh7p0aAuii7K6eeJf5qDSsDWBljV71
rjNq7e1wNlsD7c2VF173WrmCXGQEzbcTy0Kg4XYIKw5neYWvve+LWbZ5+5iBIsN4
qPxJO86hYPYo78zlC/kAu4a3yCgHPPC2BSl1qwCTmn7K73p6F7anOGaJjcF4SBib
w/XYzRxFWEWefjHNhGoB2QX5mtrfr6yHbW28Q6DDTpfS8q4Laf/v0zvCfbDRPlad
J9RAfhyf1c8yP2pIWUBnu20OUrmm5C/0MxlWhi6m+JTJoGDeWBp8KQDHcj8vYFlh
NHl71PdG1I0Q6qvYP/Sb81TjGdYOVZ/dFPcEvgDk47a8sMkE0xFtXQQix+SUSHJt
VpLJ+rsU59bmomGOZUfRVZ8TgAmgcWuTg29ADQWdilSTjChKGs0rgmpFs+z4EPT9
TOtN1qgvwi7TCsfpSstIgswRHuhp2brSjIz7u86eOUBfLWmUVw/ftiVkWTT1xAlC
p8v0iE+iAWHxriPEvmiFVhMmWFcBFT6xuc3YcC5oW35YG8LJaQi5Z4tqq+gjErWG
6Zyrm76LZcjlt4q9dRIQgW8zAG2UKEGeIjPpHn+kOp+PJ+3vzCgltZ6JekNfH0d6
UXdTJM2HC8JrSm0nxSAh34XcYcRS11BWVz6VN5OKv8wYyg+ZTs6uYC9GBi9dzamS
5Nlg64ZA7xi3RCcSKQW2EFQc2hccRqT6i4wgsNHrNrB9o6jLRTGMPJHyBmQBd6/z
L/TqrGWTDvxFxGwURyt59M2gp1fpEsTew+XfGL4H8AxkHnv/ISbSBfTHaHRggUPd
7dJpIX9pWuDiCSq+Eka7iSLzNpd0eqaFF5Q0PQrbgn05cKLnqInqe1OgSO2X2Ap1
J9UAJ0PQuWeypdA/VHdJx0Uqrqu64Ydu96aX3MonrgvkzCjHzyCyY5azY5fBXbh9
LGIrzXuJ9Ze1fXAR7kx06jBBkSc5DnCixcOJwJVMo/uR2BT/wDAlrLzTDixDVVm/
feakrJwVuq7r59qh/AODTbXdmZjaSXDth/9yM2OezCZIUlxRpgvdocHF5xnzwP/h
HSavyaSrkWhMZGicdaU/xSzvo9Wl2cOAEa+5YBoskUuDLYEBl5ut4Fc2l2L35bEy
CRf6qJBlM6VGBHJLO6xmxyQlP7jc3sgOOufsVB9H236uNa1tXk95Wd7qH+iu3nxs
62Cq3V+oTgsl3l603Tn6NRvYsQCW7vYelqhxz3Fn2Jb5H/lGVkTii0vMuRcIKcbU
Ha79PgtavDG/Qb1C2S+cTBE+wSgP0+UjQAAoKnUEf82NwORNFakjk0Sueldzjyn8
F7fZcpua1/+z8/B7Andtoq4gRLOL/QjIGjUAm0sCARZfo8fdcUl63aYPZ/+juUpp
C9PP2DQaJxOgn0PtHtrWMm1/+zslWvY2IE57opDstpJLD8Fxbk6yHiCuE5+cRUb7
178kdi4LWePbHNIzfkqlnVCWcz4qgb2yLecYhromKlrrf2d7fgZT0+GLJidPpQ1H
RgsXUiXRZ21sJpkxkGowv6axa9TVn+ve61tmSeBn1W/R+nj8luJ3m4UBBkT1lwBU
55rIXpnTe5/XJMQ+4Ru5Cofc3pCDzTrTylVxq1aFPdrtTI1VCEyN/Hx26h1PsdAL
rDdf6sRZ3UtohBtJWlVR8oDhBEtldiSue+X8ljfH2h7clOCkle5w0FZ8X4Y6t0+C
oCCMx2BVx12N1+/d3jLRZ0YqeIozPz8OUVuYMgXtbmonJPU9lpdBw55dTaJW2uhS
ZKefYwsJYMgR+0dpRf5p66dc03SNDGiMfGPh956Tlq7OszSJho6dJX0vTGxjIehw
6k3RPADQrZe0xD7suYo0bVyEzMZZeNuHv3rHspqJLdGGSnf09Qw4BGmzocJHRQKn
xB6c0O9kXNkeS2BdLqzy321omGGYlHfFseS8oqg95yCjDJeig9XuCoHLyOQj4qqR
XgVheaZHHb65zwgBdth0FjAMkqi3b9klQQtpr3rpPpOleooDeG5G4IpNKvrlwidf
cE9d/Kj7+io7m3FkjzkkVtKTPlk5wXaRsKHoCJTrXOK4fUZNLPbvs2Vrb+pX5uw/
2cILslAlAaSH0bn9xApUqminFqr/nMBrCO5Rf+p0VMSrcC1g8pdIKdWXeVTZgWnZ
qZO1Kn5mHiY1wh+MwPwfRfJjYlwPy6vdHV/6ySxIjgny9AkI/qIVWpBzwm0R4vn/
LrmhUQus3tHqmQjU1FFdrymOO65rwqPn8Jhkvq+3joY6WRSiwz9pO/+rEwaroYV3
6NiTRgSmcJAL6SSCi9icQ21r9p2ZUqUtSW4mL+9myfWyM2cSiXPKCc1cKhocKmUM
Cz9/G0CV2EYtYRRgF1Zfo5Tmcfa5if/V8MFS1ZCzXoyiNFEjPEmEaBC4gd7Kp2rT
K2lVdLK63VYsrtNbh/Xni1MG9544A3AK/75hxxob4s5dv+Rpu0m2IRR/SS7Z3MWs
zadtG7p9UdznirpEvoj9BJFvw3OiR4h8AhBnYMBCO9g+UWAz5HPyfR+L4CBxTg1A
7cdBre/rjsnlsPIsU7Ja0zL2N9/kfu0084ww6MtDVFXSXnHf7FQZn/81NALti7ZB
BnabKvgOVLGheP0mn34MvBJsGooDKNQPXG9J1JT/qoqCP1N10FFq2z4b3D25k2gK
J1GUq+YL7B6GGPZA/BlSO2moaUTmFLkyyKClLD7Pr+4Ne0lDPHzRN7oI2rD9iL/Y
Sv6G/wBoHUC8XPFTbCF1AWskmqEfXqoS0YlmTaX9XS6Jv11TdvohoyQxcqpGacQo
iHH0N8gF/NX/GlGuIQjRddneI9/bJMZ4WtQkVdmsco17HZsdbumMCcMCr/yUNQ75
HxrE99B87MKAbxX7a6iEyf6OnMTeskojL7w4RYpqX9BQhyycrRkzq0BmtiL2WGjE
aF8Yv4HSh6Yf9gIFJRslWUXIJrj3aBXMDv0b/6UGeSJwKumaSk8N24zVP0taXdnU
FUjwPmP4j/bsy3XZTvGdl6lmoXJbENZ3FewtKZRAtYW1HH+zs+KngPChvrstg+qd
RYHuBoRoES/CFr9ZFC7PAhif9oKlBXVCkpB65qawD8+Y2xTU/R6rrp1L6pGFroAH
GeRw6SyA2hlQdT+SIxqlIOu1kdgEIVpyQgfeSS3F7Z1OIH96AGvtvUEZnTZlxoEO
i8XZw5gpcQ+tCxRfgn9/Y9FxoY3hiaIHfGym1W0ZViortxf+8w6qorN4uEnxWcrr
QKPeD5CrCfqaWy4NJGr+XDjIgDZcy7kI72QAEnQ6lw/Su2Vab2EsqQ6hrrRXuVIX
IwA6fEP2pnmDg2gnlyLl0FVYz8HFOWRxtJawjzFCgTn4YKf+tB1uiVK8ykRxPFSt
kkz0IRL7jzGo0rDH4aPvtPOGtyehyxS2GPJc5rG6i2MmyC/s6P0Fc/MiNqHRpCUi
woVinJ6Xe41eoe3sdBbRBT+frW/b+LjCZR8lK833M8molTjjdD6gsy4pZKm4pfYk
l5jIs9mRtxPAGYh5RVSD/wt8tbDjoAdVBwdb0T2ex9kiiLespo8H7ul+3E52D5wx
RvU9zDG033HSwXfQwr70acpj+sSWZxExm7bRBReuGPXV2OZMukRbZ6E4Wl89sJfY
z2AL4NwWhKdD5Jq+0drBmvdUX853bajMHJ+4mqoQ9SqbBRaREqat7ZgJCe+bxaPm
Pk9IQ1hzBq5Oxj+njkT/myG0dU27QrzTSvy9MfCsbKQq+0/BL9k8k/8NEHudyUeT
tPYqDEipsXwhb2HL4U4bqa1A/NOa+hZEwX5AKRyAd0yfdl/Qyg32vv4EDwDsBC7s
zrVEBM3XOr61NWe892nSctcPBvzpg/8WqiMJyuBcLeLnN1qSLiYcVEvMlHk50wTg
1bcJZ0Jb/zil9oqg9Pkk+5y1zyb63lQLvMgd5rZesTg98ZzZfshhbPPuiIo42J5Y
rBNc2uS8PWVricTn0hJVTvgG4aO/kWZ71jmVB7uxs9/GGxw6EMoawWj8yC2yXG0o
NHM0JoE/u7KPrJPNb6ermJIUt+Oe41dNWO4AdiCf05i4Zy2aEMZzcrmFK5emWWAH
+RBg3rT95/nMUFCfW1Mpi/d6tBPIWYtMhNp0Jc2ThqGZRpMZVyFJSN0aFU0vUzJu
96x/fKfWsCk5MDYMtIC8eh+9Yx1psbKrLAejSGwcp08IYqQOQyEfB60x5aLYLPIP
Cus+IiQ2Xnxnj13xzvAssyYYwBtfydiiOQW5V9VuEaP8ofvsGOz1OLpGHQsXMfMT
r1o0oBT52sbmhBCyHXiArqC0xWGz6Ov2vJ1zKeOF1WM5E0ZDOZrYruFq5NozHOE+
R0YvkVXC7hqLDvVWZDtS0F59MQawKAsHaNIFgPUpBnIgqzdfjctoOnhB/YQ/zjMn
1WYTChZiqQjANKermZGaT9+d3IgkdBi3lXhEbPcYtwGmOn3VYmU1J0PX7hnPfSi3
D7feJOoumR4JnL5JucRCjbNaidRZ2bnLtHUv89BIz4KF9yax2Is6aU7TT6xBKLTL
SbPdJZfulUSKDm5+yMnJulv7K3zgasUsWYcLYJMY0ZRwQYbGD2a2lGgUNcmdmOpI
t2RnF6R8YVo82UYf0+PyJ9/iDbEvlz2PZwEh/fr3E3e+QYime8jxTP5lblDecH4u
bbN0wcv/A9KdLnm36GzD4hSMqx9kwEfLVPMbLCtF2ohxUcEuQ2SZCOuyksNRzRYu
BcokG4Gi7r8DeU2q6WjzdIyvt0x1spZjzGVk73h2xkch9ehxLAcgsTVFaGnJK984
wQ2znnrALe7t8SNsGgcjXo55HKAJZv6mDJuBnLywTbAEMHu5+JGQeS8pc12AZ2pK
8DbpgBRjuVSp3dxPv91zPg+G5SDtfN3FkLM1B1HXGu0e+tvmFTb2Axx/lfNVIebM
+fXreJMd+XhFoafZ0yllXR9hGWbQOsN7bbVsD1334sHcgahzZTg86ds8mKpOFh13
OXE7jsM81bF88+fBog0REtVngnbsrSXY3hMO/Wioe/7amh+nX6SQ37wCa+gt8dht
cxn9r97YSvCOstPefttkx5J5/8Dyt7vG6K2saF6WJcfOh+r1cSo2LPSZD5myimUY
D91H7HwndcHEdw+qM2XBaU6bQLZ02CFhihwNrnFCC0ei6qZA9myrn4Lvnq93k1/V
m//MLFEaAUxgSL0ABClZXB7NG8MQFV6Hcu8nepKj2dNpkUNW5gl4Ub8C/+tcdz3o
FAThBVYi/vewbX1b2q3VcKhdAYxs74enLmT7W4aJ2hCBy6q4eCCq75B7F4qpEL59
ET7mEPXaaCJVW+z92yOgwlMX+YCUIHDCjjfD914ASpQuDyE5XoHaKTfCsMtBQ/55
FaWKoFygUTRzC0abljJhQW6+nnwHUPhsUr8lt2eKBVhcq14DJbzCvxz0bcSxzQmt
w+h9hjZGEDMlhJ4ovMRFlW2JpPITW0WSkd5p5GJDVRDEknDZy8Ojz/q4/Fxjn40k
vHFMyzoGkqA6kkqhV7qIDwYJD2W6ITbpkGuqIR7a6/6XA7vXy+7pF+rLmEHvYFoc
JflscdmKO/rohsdZCODn2zEb8TkRY94Qh2iIQgD6U1E8iGtAHsxT7vK8eeO+cDth
MjebEPobMOPeUU6EAp9XirGmi6+3oTHC/kbclgauaMvlK+3AWC8/bRfdaPmeJe73
y+LAkSg+fbll+aeuoNjiD5NF5Ad3cS9PzAwMkwzve4fWS1xZ1XxfXzbfcQKbGbi+
T/K+eDH8rX2dEnHAeA/jEuhf1yzdAkEo+soY6339Vvnz9o17urbMtwRv+XQcwrrG
ySk0EKUmxwME5m+nDbteh+9jFGXooANg56Tfl7UuzuSRdy1BFeEfdpr3bKBR3W8x
HSc+fX9PkXTxeFHKlPqNd3KEhR0VWNRQxRPQDq+Ke5kNBMhrfGYl3RvjeTOCy8sL
kxpI2rVnJzCKEs1uDNQ3MeSYtlZJXNnIIsf5NPZiZ1jmVhMx2Piy0M+2ZHpPQ3w+
DyRChbXsl9ga0UwIRVH6weqcQf6mYXxxcljzrPFu94H5K6uXKwsFuCwUWREaUWfr
OTIGRc5nBQ5Bky+e2K46Af9AgZ5usaS9IX4+TNmd9/YSbYqN25pcVAj1LfLoY1TV
JmK18hyDDjy21Bg07QGg8CHFpGetd7YbC7gZnC9s/POVaGs0tslQa64Vb4NGjvHs
3V67Kou4OXdvDCLKYmlTPAcpJaDX0uR8LI0PEHz+9GhXGHrNddcPo+NGPyOApR4V
Nzsw1g9yto2+q8Y+f8p8FaNZSuossqIKEBOVJQtHinEULrbLZGLkZNHsbb9TwIxA
D1TFYiexJlRRU17zAkBWaV4PNFJRZtldIWzDE3V0ncAFsp9C1hG3hAfWQaZFGC2q
xYC6e/ouzkTyH+uwuzrS/O/lUynh7d2WdMj9R/MJYiJ76V9XKIq5Yw1vmNZpitaH
TYgtKaUAnqW2i47/bK/qyQM3vAEcC87M5RRTb+22F4Unq9KCk5pp2sJ3Ncu9LAfj
wRBsR7qY162BU+oXw9fhyg2cCc6PTBa4ryNeEgKaKtr0hJGDaavkbhbB6rP9Nj49
SWG/pNTqzXm9v3c5M7J1rUHhlyzeaFlK1M6F5KllSLnhVez1ZNqw5bIb+Kz8BLTJ
WkGM9dkBlDa0bQgtuc41RqbeVOzr3NSDLhwe3CV7i4IpuGYjaWMn1e5oaDX0Ogin
6dY3rYhkqCwb2YKmpwkQPN9sVyLwnIK3to64ExBQvo5zau2plRazqTA855XrrtFG
QS8jad+ysG5T2y2/KVKgMdtL0Gi36CTI2EojwNaDD0Jrszd9+8OYI9CMtTNVcv1H
fEPB3lrR6nddILlKvjb6j/8MMq7Ma8vW/03A+KswvtXCXqQlNaJDyQc5WzaXSVZa
gKVPLb8+NDU3OaU2uZh1v4OHZhLwK/YbP7eb5F61LnDS+uVaJystst9G6rs1MAGg
LITWir3V8NTH3AsO8MSNwesi18osiccIzrzzIRLh39IqxsNrWpqjQcqah80JBrcq
KCG1lLCEXiSc3SVYnpLpdMjiiFY9+pIEdCSYUM32e4P9YLoxX+Oq+JrOb74PPw4q
id4fJMFx9W2wBCXvaxYZ1fxgsdoh4FXeIb7Y7IYAS7AS6I+2fVrVzOe3XO5vfv4b
wTWAD+GUWgGX9sXj4z32+jTykNInc+D9gymu0a5uCngTBw4lhsgP3p22QQQPUnuo
iHTrzu9ecGWNplSUKyI50j2W+mux4hN4waasdgwZQ9zPbx1S2a6nmxXzRRUA8l5/
B3FaHII7F9ciixg/wXSmCGsBJ881GwbakS7hfFLycfZkp8LZIsCiQVZu64b8VRxI
kfe18tU1TPV9zsNNIAhUDmyQvi1kNB8Q3HOWQ6udyvHCBiB92RBpiMejhqcIwt0v
BLXZv+TpP6KkTW3cT7hNdZ65lbgw8t+8QLQHAS67bxpdITJxzI/AndG1o6LkJhMS
CJPv1MwEm0N8s6a8hG5gSPuOPAQVpfFz4cqbMbA6ff3Mje7aO/WZu+5t+cCrfaRz
9ljAp9/vzh0H0dQl+NzEsgEE8rEt52wGR07xFCFhXkT4DMAZSw5MoIiPOQXgrIxU
sI7C7pHB+s+yQXAcuUYhZdnxxrkm3/NmkWapLw2KCwK2CKSV99i5C0y3sa5pkg/c
0/2/uoNjEPpJczasSHVGIJTxWCGvxJcwcP+cOeXeDH9yyUwDOxzwZEb+ItoO22mR
FNgH82emEawbiRNg+TWSKCiMvepbkLddyNHQiKpL8QvqDxx/fagexlse80KZFKLc
6aNXZjQAl2ZkX1XrU7dzUAnlRTVUhdp9WnzUrVyfxsLxjQStqfX5QxpwOZ1vrTIu
HHhwht6D325G4QbTFIX82JVB4vxtHr8qRsBEwWFQvmxRLE+QL2wgupLchm5Nud0C
qI2G4OXRaCUGIWXd/7pu+MkWPHqiHPwftpkiwAG/zVF8e6XWoc07uftTgkGYxFQV
RkUA1EYKIJ+Z4ZMW8A7CpTiVbD5Exiy8mA8U9GpsDeFh+LzBylJadc7Ev1BlX4GK
dy9s27uCqkepghrpUP6LfM7ltX0MzDXHO6WjR1dwDk0bKlNN4BJFljeAaameLa+2
eXbQlcVh20MIzLgGxFAARItiyiQAvbRJCFizEyRZxG94pPHYZe8VagoHecHsN9a6
mgBpRqWuhGiOqQhkG9DD5j7/x7S0tZhNKmb1+iGBwOBJOEq0DvoUz8xCTcCRUVRo
1Ca9tQoNBIdd2drP0YC3BHYpLXcbvojQO7yDAmjdtXjQPzXzGKoNNc5epYEbX4Oh
koEax5F80Bd4NdjTuIkNAjkkfInNYbBa2+bp6nrmzIzMLJRhel4VWxqkWpU1/AXQ
U2bSs0BqtAyMPnFpKcTYdiSkpR9v6k6EhGQP4RHcCwqdNu9UBzBhkvUVmW/ZHWI3
jbVcJ4Ug+Nb011ap7sIJ4q5ILOiK69x15USyyKQ2uicgH9yi1gM1wkGSdSp/N+RP
Y8Uj3IA5RhYvUK9woykzqlXmqNe4xsbkUphVL88JZCWH9dwn6v1oQBXjN6lvkt7c
vtGAu8fR2o3Da/zLPp1gyQ1SQ8NwLw0haPpCNRt/x4Ay4fdQ4A0jMZ4joqyA/DSN
rvQE7ox1psq8XvU5jgEDvA+JLE7OGJCVTYxZn+3nbcT98HclWpmRFh5uE3qEZol7
Uw1RDAadFFQuvivgirrEr3dvlcA+Ro/5Gd5C2dxzX56VWOy/a5435R7WzVbXNpkk
EXV9Hiku1uNWC5hxJx1WBAMAo3MJTTXTd8RadvgpGj6BSuhjRKy1Nk56gVjVM1aM
ajVw/KcO7J2kbOS2ivo3Zu+1Myh5S8DzcTpGJc1F80fmv8NXkml5w14JkbxUUNaX
FaL3trfLzHgin4s50FPU+yxdNObrHY3GmO9rdNtwH9kl6OrwoGrEcTQozzDtKFs2
ms8oRzR8287RlHRvbNzY7gXQhGe/twjwDroA5Z4+mWFzLw33b/adEPz7FnA3prpR
xgjefHsC4EF8JEDTeTgaKOfPwCJ/hTFfi/iBsV0C0W7C2ijjQKi8KtOmajdovJ2o
cFXPOjNQeCi39iZnXigVRgY6AFhd/E+MByskeZldhurEGrHU6H52kYnHwQODSUgn
FkTTJ+S3ZytT+/z73erIIIcvu//lMjtYq30CLqpO9zSc1S2jD6abwrBLiZRbQdr+
KG0x4UvhInOG0MPCNACpZvG0qomA4OF9ZKJ7mPLQC8k+IsDkRoXhSGk/yVyfrY1x
toHs48RyLMxRdgpUwb/fDonwfYjfjCaVlMNe9P+HCAAhY3/bwSmVTMOLuWdM0Av4
ALPfO8xOELItfZ5BK5Co048K9TCFeITfWaYnOoMlsKoyTDWwpWB2p8Dup82jV4Jn
kklFjIRZVjWNS7rfMQIghUMd4pdfLEOKXIFfNaiXXCRKYI1lNqyaS7riyOSpUopC
rqUQtejUajcd1x4kpERYswUSjBdBDAV9ihR49AAH29gvU69BGtF96D2LnhSEb86I
tpBixiZxToahqlcOmZ6wSSKRbTwp+mZndM9WpauY4/8GMJUDQ3OAPdpnB8oYq5tF
o76Q4cC7vJpnVPrH6ONPulR33si/YwGqp+8O5DBy7uc+FPHNP/vmA74Rc7y505gJ
orZVWGiAX6y1D0J86Oy0DYAmgXOuDluqhxxzfN0Gzb/VA8lafobjJpo+JOWpnR8O
d7/x12v8B2kse4ox9VtnGv+Z89exW44jwkfhvU2QglKjetK+2q/hS7EsLOCn7Lqg
UsoFRx0TggqVliJTijkhvUg01MASyIIjHwjTKicw/NyANoBoGjp+9XW7V1uFi0mn
yOQRsDmJJak5uAbxuwELkJwvNYUUu9kQcS0UQtJz9Uuze43R5C24G/JXXb+Df2e4
Ilf2j2WZrvn3+6GbvSgZ1L4rmaIIq9c1VqrqF7ym/sPhuDakrAHfPEn7D6prbe5r
4AwfYm3dAq5i4gfkJLjKs6U+6W0ZcZRsFQ4i0SQLUIckmNgUXjBzSBdLzd0MlnTI
VM80nfPkh1Qqa23oPgOQKmON74w38qbaVUNRZWw5rbd3DuG8ujruWKdSi4M05tJG
6x+3lJgmbBRDMv49behFRT21mdLjFoiQUC8NC6Oiw4aZFDh6dkeTz8h7nsMtmwIL
SyheX2fTQNGw/xNcARPtiKSc4agkSKxDoxLjUdMmcnnPAIXKwXi0EKVpckn5zpsy
SpHdx+L//s3i4D8XyKrC9/nIppWZHoEugph1HcMaMLpAMk+9XnAd8H0CVOBaKN6x
Oq3yPfoTc5RAiEN3zfiAl9Y0krFBaL1IPCUZcNfp/Q8z32sQJF+ZVvvDptw6vZi+
zG4VWvzbUfBP7mmBJJVpCtbKjXd4NFu+6f1s3snxtLAdjyR3b11qEf7nMiM9Xr3j
Nrqjlv6j+FxzBQGobBdtHsP6kUVX/IV6lLy4FpaV+pAhTn87H7KTZBB9yxOKkMDy
B91nTc0mcADgSoVNPgPtSbVojmH1nEWZYU/3RJVrsXkdRTIvTS6yloyCLW5hqqSy
IInaGgBegamgoH6YImLrhtrCqWByNIQBMk3EYeEcPDn7B0/RCN23yrns+B9NzhJn
pjfTsRzU6FlovUWQyL8gnaO9Tud6fkNUfEG5nR3w+kkpga9wZt0Mlrk+jLdUtXEK
6VFjk4JOKuXumiOs+iXkEu/DeIv1Vk5Y4gS2UFLBvtLsiTQ/MoeVs8PpUgbB+HXi
Sb56WIU5sfCcOO1BkPXlLQytYfZ+hYfqGrvNUJOSQcAoPk6zTj0f8Np+4hKvvtnH
/5iTf/Vwq7YKuKcww4JVcBCYuFIy9sLngCQ8elYYATBeVzq5+ihuAM/JrDXbyGxg
JbWMCcS5B0oafYMeJtbTv6jUusxZCkjwYm2Xz9mz9TcYgtBHj479r9TvlrPTwPua
j7nrgKnue3mjLoPwR/J3XdY6CqoQft9ol4SF0zUTg902DibywMIV//pPpjLo1DAi
KVIvCLGB/W/PiXNW44YFXhKDGEwDg9vPSjp+ULwRGp7oTXF9ZyAkhQykyIQQtPsc
pFquDnn2ScZJcQRIqMF2XNp4p/4FeJ5flhF2+LmjF+v0l5r1PnpyiRxC+riym+MK
v8oXuTOa/U0SYxBPm4bAjiAag0SlD1cl0LPZb09ScTxLS04yqKVA4GZBmmD50Mqw
RrOwSQu6W5UynQ41H/G9B8v8d2Qokh9aND+h1J1QbwSIu8tqACVESU+Clj0BSztY
M0wC4xHrHLyQV29/BjLPnDka76d0XGOkkLXV86v/sbFHCw1Z4OSEyDa9EHsXA+s+
Plt/lFdLVpANlvxmsG6jCO+wj25xTDDN2RARqoAEijZe0GKGrEkw63B+TjU961jj
sXkaVjQ4RJnQ/L7NaJn5Pq9JQ7QMm1tyyXOVgepywY2T+tBJZF94h2tPFxqd83ul
vNV2x/vnjOfOjXa4WTXFZTfZ0XRqAOVpZmZ8Qk0rgk5OQnYESsa+QjLJdPA9CGCN
7mhRn/s8dUWf0H1I5HZV50Ndc4v2JvDp1jcqOmtYBnuioEmMNni/d2uJBSbJUdK2
uyUkg5OgNDuGo0mkAWe9LyHkBis+gogARJnvbBNjpk0L/Pto87bn7AZT0g7MdOq9
mYDjNAmdNu4TaSwhVSw99XbCHxSKVNgM8dIR1Yh7VmoX3DMq4Z3dYEmvXnuVgsLt
96wpQm3mjmduFOhkMNc8xRrKt8VTtu2Oxx9NuuOrpxCjeNJDuX3I3J5O0ByFx0Ie
IVkWE8lXWWc1jd9a3/zwdRknAMe0HzRnPy0Yt9rLsikqtAbbN+xHzYdiJFM7rKEl
+AXWKeAjQqHwp9p+ixeTfwPCax4wsV6XuY9O3tTjwfO2ivWEPBrUhUl0q8/Zf/D+
+bRpzqRvV9fYTu2gF9CGwVmBfTPIzlY2OmKrpzMvIU0YPmoRrcY+rTwsPMsD4cJs
wEnIGaVYmvvg2/A81594iEPKdHBf51slP9Oo3VwxVge7F4hXtAgHPh9VrwFhfqTJ
Vo9o506yJbjTDAnBNeJU97Ic/zbYD+JG4o/KCw/h8GvUKCRcL0QH8v/548balnqL
fsYGOwpz4KeD+NaBOz+WC96U44NL+oxuVpjZnTSEY5gWTOQ/4s7YqdYJSFuTiVoA
W9mr7cZDzX6vq+WHazMDoFNFWQ0lDUGMlLYNVIlUqLn1fj69fbBhQWNrkDkob2Sb
auomMArKiOcgd/96j4Yo9Vb+oUo5wvHqhFk100vAeIaCtTFbLUoOh0JT9ef9v1BK
T6TifvE6EeqqaM2ZI6rSbzU3SvhlGENYgRLLQw0HGh4gW1sZeoc7X/Mo0BmejN9J
3S4CCkUHyA78iEFFrMugWUktydZUHre0hr5W5CrMjuCoFz5ZFQ/bh6oXwrty4We8
xd5RY+2FbDsNWvu2s7BUsGQegGqa05bY9J60xXdwTkTtc2NqIg3ic4nO36dCqeQR
EoPBAdqJG4WXmU0GooqLKCXIw9EDcV8PUP/x2nFWuZejzl9Pv18zDxBJALOVwZU3
H36gjvY2LywFr9+Dx3ElYTlnDBW5G22y1giiRS1vc+6LFl5wBl7ru3MbLlrZqJBv
05ydzLKNBqxzSPlTj6N4uYyJcp57r+ECk2vs3aJbioOnMGhPQkO9l1apo67qmQr4
Bdc1jcJ98neLIAXFch1ioBH0RNiqCC4ZfZWzKkf9WL3cMXjqe/AJ7b2dAQzrI1oI
6CSz8HgFC3EIakI+U+8JpGjx4870sLGRz/AJFeaGKIduhHk9oxXnAeM/UInA+79Q
paIfo3ZJ26u249J1fqlJDrlMhv2FMb/ZTOHAX2K/zuM2kfjW4hMAjodYZCVuewnK
Z+5yqiqy4RQD1kjTrBULcez9e8TQct1G2qh8pl9loDoS+knl1L3qCo+e4r5TL+K0
q1rva+c7S+RyDhGDvnSDtQFzW00Amenrw/1y1VuXBejro9jKau36L2HXRXv54DJC
MfR/cr8jc+AIW7xXbCRg4SHHj1duIIl/dWYcYOadrlqXpYx5J1JYs4t3Q3bzjnd9
hYSGdbki0KNeeThtZSJ1iKP/+THXZqg8l0HkCJoGB0Rf+08KlkexNe/Dif7rI0Lv
5ILx3SXku2uGTbng8501DgsxMjSl1iEg/v0K77BbnaZFEPbvOSucqY9PfZDbOS0J
6LGjS/Hec3gwXFaLkCPFQbk114hME+adjPiXxBBDJBqKjjJBy11yplI1izEzydN6
e4xgMJ0PXPZDj6q95ic2H2EvargCiY9rsA0o2pPo7sZUNRpyplzO/MTuvD72eE7u
SZQyR27qbuQiG2anRVtZ8XXjzAQeivFJxFX5vS4M/mVkkgOhgN5gOkJQzxdZU4j2
hGLbLXDyBc+boBPKrtqRju7R+MNRKtgkxlc9ksKyo1G2l8O601z9ZcfGfJSpqaqU
kfuQqlssJPrVAWPfQ7srXTMKMCuVZmUu7x70P3jmKNLA58wM7nz9t2pVAIU1OMVL
o0w1HkhRpOSPaJilMYIBPdbN+LY1CwvXW/kOKcWEoGBd3S2OdJQcxyQ4X8YXjom4
5xAeJSBHEBw5acaByrdiwn1bF0KSlEIWOZsje40V1flgnTZo6ouzdTezMFTp35E8
hyx5gEOgT5GCRpke7uMryGV8Iwi9bOFou3C6J3V5YE8+QjtVk0c6/uePPKzF7Eo4
PUxO88jTMsU9MyOad0H0/eHh4u5HkLr34p+e1DHgeYIhJuGrP6viiBagV9MlOC30
fqewRGfA3i5QloDQo96CenJxPxDXiXMaPShEi96XJgeedEc8D1orORUWWXkaNcIf
LaPyHf8rUdmvUmCRyea5+98fp8mU2ULEZDRVBtEQi2lix7bDTII5gGirHlrv4IRr
pX7A5DW7ckhRaUubK21cEyfi8sVf0reqh4oFEk3wNi0w/qtlPliIxzGrZa11EWiB
JwzQKPVhGjkE/vFjJL+++x7fmjX15zy0zzcIs+eQ/VLHhCj/Br6aP98GoIQiHsHZ
ot3qY18hD5riXhkpsZc2qvp/5Z6jaEehr95INf0aQZwl/HSLWKllJqRp0kTKe+Xs
hZiR4rc9V83c4nT4Mpajl+XS6ZpzNpnYMzTTh1/0Yoy4dyxdsYRCAkfNGU7FRvp3
hTUL7+540hm2UeU212kSQcZf10wr289JtXi6s0cya1CVr0YkSs7jIiFlbNEwUQkt
4WtNpNkR0zPqUtsYhK75kuReuFSE9KjKbzEdY5T45FzEMe1FQUbEL0ftq8ksopfL
yZGUAnJHwqeMHKwQYJqDFGhhWHt1WzLAtQzPnJuRt2ZS3z3SAQ8O9htsXNFtXm9b
4rE3XyTXtKHQPvF3ExR43HMpgGlcZxRpW8y00gWZvib9mS4zAOKLeznmHetWIvS4
Vg+gPe6aB1uF7TaQPmCABNrQMIwH5KinxUtLpZL0QoJr2W4k4VIWotpbvZVB5MNW
3fQIcydw0uzHOkcdQTLbq60wHPLKFPfAhjFNWHaB1H+FHPKvBlnDPdERtscoIXzc
TxJg5AkdzhbjqfmucPGnnfPij4FmZYW8Axwc7JWYPuR18sv2fD8lgedcoGZImtOy
F1wMfF8kv/aHXLqpKsibHn4Jyvf2rH4CvsflgUfODaiiiJtxfNanpGiTB09VLtDn
EVr2uZUd59C/TSqDPNcPzFpQS0gLhFCPkkS73VaM02qASl+rb4gKgMsE4P0kGDt2
fPWGXDxxg81rInoGTqGB7tYFyo72PQCB4HC0h7NLulAN9d8o9/Tk/O+Tx2/YRPzM
7NZy8QgxTvrN028ymePnm1t5yMjqVjUCig7r51bVQKdKBluXoPhcymrm43PArvLC
P2ucjlhOU96kLd9jJK5Ez+ZylxfKxF3gEjVC7pn/rtIDlzylKdElMJFFe1qOjxaR
O3SyHnRKoS7ul0P/K1Qe8/QVC4VeONqHNRyJFX510M1gzdJ4Uv8IBCnd0ExVDzJ/
YpUair8lo1SveYI8aMOQUlrsLl6sD+K3RQAQw8cgf+dPvawm8bS5k0eNebIGOd0f
dQ524fxuyurF+vERjiY2YILjGtDukJ6EBtRnGjwqarVOCCXKDIvGMOLfGbbKgIAb
ofmQNLd8hQ0+wGHthOCkadgU38fZEqEff2SjMPQ03Z74tTTaxZ8EsjthC4e8taC0
E+c5JOtF+RIkveC0FI8iVc+jX4m5n2tK3bW5OVJ4tC6INo1i6YuIksEPg37pynjG
XaQVIAQGYRGqC4Fc90Ov5BwXZqDdeblM1CNWeWWLUmPxugBXWZpa3uxuq/NpyFtj
HNRwLt/J/jNR8Fenk6YLL2irE4f7gF7JFR6DYe9cO/2oxZF/50YJ+AtTTEMFPTHX
bkjs6VDWdwPVhFDZLTz2bxQT2BAbPNWvSAJlBy0x/624juiWPWf2XyWyNTNwea6T
YMrCGSRy9y6QYRfHQzd8kwXqcw08oBY714meqhG/Y3inc8LsQnr/ShdhrSE6Vae0
eBwo4SgTFtA+NPRzFef0lxv6p9P5ysyDDrr4pJ/F4VmqUgF160TGJhL/phRoklhS
M8ZQ3oWNYZM1lWGnwl802oQZamW7Nx7aSOteXgxBaYvgdV7ewsZFqCedvPFI7Fxj
KJrSBpOhdukzmyzf3bkzwHk5y89XYy1zRGhfIjK3eEhk5wzh0tI0k3hbb97T5xYE
Sdbu1zNhHCs4VdNizAz9Tm8Tvubi5RfsULIpWOKMms+95l2NFCoyJjKU29CMO6Uq
ioTV4ZBkI+o1RBizJivUDFyKvdmEDkPBso9HwTdGxX3jWkSfyinoBF2GCbeza+DZ
7Ni/xlFMLHh6rOdJ3wVMpmVfmAPC43dt0lhMzkqzbOpe6TAPg8DriyFqqiBM0WIp
zH1qQU7GNUfDCL5zedyBRiJIZ6+pbgGde/NdYb8niW10k3lw05InufFuy51svZt4
Vkr9XqxQ9p12WWfKwcGl2XcB5qUCdQdlHc3dCitJxAjUylJ3SmJfesEqNG+Q/9xM
MRG7KAE/lPntBVLnrzH2KfcTrl+vc96e1ux2bxcVp38wUoz5N4VChrlGXBR8Lufe
v2DAJaw3js46TWCsNpnlkZ2/KGB1lqrsiBRnKtGmKFwlrC+eM6j6r1ZB8Jrxq7Rk
UXC+snoTfAdyz2MjC9zIVX2W8qCrdsczRPvfA+F4IsODziYsvmzOGTIUx9y0Uqpf
b70Yn96B3xs33t4gviigb2UnIK+WF0IkfHLX/aoE/WVoYlZ097eNgHUl0cyTujKb
cDxt5aUXA8HXyTmh8da/6KfaStLDlIpjnFCABSD5DJaMbM9tXNf3Ohk5pUAi1NE7
aAid7OYwdNuAetr/OPZordWBooYeAqElnTMZESI+m4eaDaWfafcYNbIiw2XQ6PK1
X9e+AB7lUE2XkILPtd20FnoC4LK8Mey5awsTAIPpwtLo4kNqyqQ/70o/QGR5tdoH
m1zkfD6HbOR+VU2Pt38mkDmUgDVDe8C5HaHbd235ujLH1fjCpWn0zinURRmwccTo
PZrHn20NgruK9zQkSASvq258SmAdm3RVE1zegfpt8fBmX+7U58JI0w+o9fyt6k/8
uE9jrQ7DZG5whxxD+gK/eFK4dfEtGsGx4lwOTmwBZ/R2BhJnBoPXKC3bQhyhgSHM
5y4buN7yZmVlIA7IQDdbz+asAb2GL3WVbP5fghRs0RoHjf3IKZdfhZkvBVCmExa6
gPOvOIcU5PLWPJdZpWrjrkF9urdUfKcai+bO5gZbdlO965/2p7NrRpydvWxV2U4j
BJJuFwv39JOJkBDxIpLyEsvjuXsBS2qePENV5syDpuqxdlbk9fuo4vRs9LQq1/bh
cSP+CTqjCwAroG7/lPv3zcyEPF+NOiNjkhtgFfVy1PHKyIz1f7pn97GKn29FSOEv
l0LyJFfXh8NO69JK+n7fsNdNuTFCquHlNfkH2I7ZMIHbImyGvhnty086ArTOg6gA
d+Opg7YsHPumICoEBsY2l66sVPYXz9xdkDeIu/zwkhBSHtRujR4LwnyPIp2v0R84
YycPZ3+seRNsOjz9vwSsJlkQfv1EGNoa8PkjoNm+DqnagI7D8P9M+T/zLSKJvpcp
8A7ouHpEXXKm60RNGlboX6Cm24P28+1w3ODQV0Irpk5UmHorsvNzhUwiMohvp63v
kqFvwJ6VBB2DyWGvl6LelbyhtUqo9qN+PqN1P1mfZ2KzWxC6cw3rJNcPsXuRKgrH
0wO63m+Y+YqSkXxw+lx4kkQGJMj6k1thLc73WTW4pC4FeFN6JbLmadgRLVKekTdc
pVQPbKGZQuGGwWQakBzXSspLa5YU+HpZTiYBY0l/8xTDp2XayYYtKuFgaxDWT44E
LL9Wufm2bWkAlY3qj/moozAZb61SRkgyxyjkwwX8j+fZz8SZcbhklTM+5D/zkeos
o8CCOTsJNSGFvwiMbNdqOyg4CaQNR8JY/q3h30mIB3jm+r5ixCFwUcQ2tc85n/7p
eHFPcWp4GOcfmmoLTgo98ueWRYQfNGXr+gTSqb367BJgCdDcTSJM3H9wZ57LgQiP
wEkWXnjOnW4k4/42/AP8VP737v02K60H6BBhToB7yWoanBeuKEVaQct7XafERqsb
DF4i94XUqOJjJQpvBo0lhA9X3PI1SRzQ5Uy08XDymWeGJj8Sz1Iw4BqJ0Qgxk3/M
zZwUFzCN8ieLKyKwA6EYBBMyPAVapwHt38HfxwedmP7NvxkJRD9NEKUYiGPZ9mgx
RohnQtjaMdztL6E1FIC/XufLikKAyfUpkcZzzRnCX4Gc3bNROv6Mu0BuS73ST1WQ
+Y/ioIPXOphXeVyXn1Mn2LNdt1hdTd/vdEX5y7pBJYdMH6KsiG3z0Bz2+cTLEZSn
a6J+R3OIX5chAVAXrU7ToXSFWOEx0Xd35QkIV7qb7cXVKeEMVLd4Y6OAJKFVVk7u
lxn2Y4btAxkHc2s9MBHK61DB/V3lr24/hWx7pcDrkKmIbo4cLv0hVTt+bMDLm/0z
ZVBmjWB7IAp17tt3a4bldLrj6GYFNKz7zJS1zqTArt537jP0Dw96vir6cayErRw3
qqChZNKYkJZ9o/dfFrFpMJcLf7hGiPPvVYF1V64suT2PVXFaRuKFzojHx8oxFDAi
iEFY5AfMnEPz+dR4WUP8Ke3cvd3ukoN2smzrG2UtjPjBC6GNdtTCl0iC1Ar2MCRc
devJjdPXx2Ec1uDfLkk3Cwz2ug7NNroRevXwUAewUnH5kiSCxfUBmxyl9F+WV715
9IpwZW8YhZyyuEdmvLnsDJ+JABsq/9Z8qanA/VbtnAzBO3ab0BT626OA8U9Pvn0+
jrGC1N+nBFyWH/7asmCyEftIA+jH23Wo8twJpdsJghaO13DGIbECI88KxjqqfLQs
sNbVUtqJrvv/w4rYmx3BaG845kCdTpFVniX0woj8nsi6KK9FEKicI9+do4EBOIAc
GWMafOrAW/S3A69J/185r+E/buevkYYFpViQPCyf6vfE8zWn34xLCWrImtPTCnq0
/5w3rQIe2j50Bfk7hcl4RMRN2m61kxNA6tn+mSDeO5s9ipM6i6iw+OBsYQX9JLar
ehM7W2SK18b5OS1+U+xyj5OYojnSCGAKeujPDFwLi5aBdFq/xvNSTamuZrwNcBbL
erm9byZ4iCEX/mPnZ4qeT0Q3h3WNchoD1JOjM6j9F0lljc5Gv0BNXld4EYB7y0Di
s/Zt/M4y3EOMGSbvbsDAFSDqoy3AQn9LElg1kjTaq5x9RURSODBZvCS6xJWwNAJy
KhwjWw/KMMxDcwknk2vc48yKNhgMZIUli7W1Ay4yycVWU5/wSgFcZI8XgpYaggSy
HD0WTHUuIBEiZSmvj/TVy3MJbzu1gyJb8z5qtjDHhznoo8uVH/GoBPtdRE7gbIH1
j7o2DpRTm0VQRzE+CkRG6SiVZ/73+H6BkZUEd/WhoPXzSpVRq1SxVnnx0E6CsQOp
xEz6VQHfjmSukndq77F4BbHNoYmRnMQ5lseFO5se0LuDBT7h29cd6KC0sL1+xdvo
85tw3vF01X6XmLfMHZUF2KyIorgi+3z/85mayEUWvr8iZjGs72dmpEsEHN3/paaK
S7dgYPXGkl0N6D1XvJmaD1g3JMzWAjVhuiuELjPpj+6zd4CXS3sSFT0/aTs547lM
9MtSlzjYZMNB3yTe12tpFMJbOXwRAgLP/ObnuNYiX08T0FSGA6IyjiHZ3Vw0wNo/
czsag5MDnSGl+j0V6dTp5hD6jdDN3bGH+W9/zxN6cO4cj/QpP+gwwfkHvh43Y28g
nfCbywj6Bn9b1lqu4awdE9CUCm/U8is5wG1jLxJmOys1PlsfwxvSTUuyvD6H0yjI
kvMxJPmM+6JittnxSd460e390h1IMB0eteyA/wZ1TcFpRv/mAk5mODNcoOLALsz8
H0vItzR8S/M/fkuEX8yb9/XznGxzxAFemZVep8MWfWmXRtqoZh2WQd6bUbLQfX/S
Ejx+BHmAnN8jM+DzlTepl9DPF7Fis5xroAB8NFSFKqIcbRaSSUmOjhuD13yvb62N
2NjDFqZeVCW2JN/33nbzKepl2aaNO6zHOR2D/nMWX2OVSqOfeeReP6wkVQKSgK/I
/ICYl0TYsZHSB62eWfIZ3bWxJvO3nF5DPk17wBFA3Ot7UQtGnr5aM5/YJhDwSdvM
4XzTWNo6Sr34fiZn2BnnWZJhp/j6QgZoO/6v30+pzDKERz00WY8ah3HAUm0TUw3o
ReUyoevlFgwGFY9MA8njdqZqYjMXxt92TqeUVWDpeNzg4spaWmAoF+RWIffXqQGH
RVj+J+rdRC37uNBVi/Dfu7XedfcDlYJVHY7RQXFJlucGGIJZcJ93Y4GwYaw2ON7c
E/4PUNsAFg7It1ni3TCN6Nfomyp8gOB6jFtA54DrMhDGWLX9AxOP3imSB0xIHHy+
xrjznF6I8zHTI8oAjLSyT+OACq5WW8Ek7jDwpuLdLgvambJMW3GF9Rffz3dtQGpb
pdJTctXJ35pUEbj9pmhvu29PGEtuKY2QwlLbromJJWGQ5dy9r2VZhn6yjHgZsoyI
2ywCBmnsIg3hkREa/3dKmM9f8tQsKTpxb9vfgI4sSM7Lb1gtp2gtHnHuTY/dGWxI
oHIA9u4c2iyLrSiwah+qsUTwbyAz8F3ueVqu9XY8dpeYAacU22HBSEHAvXSDP57Q
x3vyM1eOIXGPqU1VtzrcgJy0v4fj+UucRUxIqNyp4efYjtMPR3u8W/NL4222Kte5
czlfO5KlsOQ1TgzYiFjohH81IW+dp3fo7tAn7HBDnPumE8QWg/z4qCE2ejVoOnKM
/m9Yfc2nVima2EI8RHS2r05goH+8+ZHX5pjNXriz9Ukvpi5ksq5kHbIOPgDv6rGR
57SCJScGeCWzGyRCUT/GOxbRtpdnlfdZbnEYD81TG+N/2LngD3wAdXsnIlL3HJKJ
dFCiUu5occ8Gwiqrj+zb4OakeAxAj1l0JHselUmhAuN3BIhVobID8dVAhh5OAeaO
NszU0RgwKEe0mpOZdskpH0KNFY0KGEGr8Se5zRZ354ZxA8lZqK2cZQGle+UH8Crp
Nc7QaGZU/jw6zMjh+OGXMxtOVqfHmxZf3PTLFLFf8rBcNhmftWeJB3XAywoz0n2T
1Rr1fm/SZ9gKjcd6XdKje4gpE5Sk04hSBmGxMRjIHuTZyAJEWfmxXKZfx1oj13FM
Q7+qA1SYj/hlS9FLo+Eq3sHuf2YXKls/5zE3sL+WxA4PEgldmivJ1/45pxLSXq8i
JOo2N3hUMmyuGEVnLZbcFArq25dtCOl9JrKJiNDXoOpjdrh6256MNKHiL9JOLyz5
4fqSQPHZYKBqMBYN61BYs9Cq6p+Gdh5m/yA747zIQOkPaJLwiZ/8fzNveuy74six
WCKIYDapse9B/rRSwommAkOPHuyytgI0FpIC8jkGW2rAtSwi/f/tuxRIoijuvdlq
UsuXMtobcY6WfVa65TRG+JS953KayABvRhjUQYNq0HDPYtJ17MD3jjAz6586YzXo
uR7mCWSMm4nfjALG17nVmFBsXqXzxgXsUKWOcFnrnDm2AfIy8MFL5U6aWFkg1kXM
R8lXjxtitDv6V7egOqNjOS8NIKqcYPgqlI53VjZ/n08r4A96qstrTC9D3GyWykG/
lhQb0p5DzBs4LQksKY311yczqjFWKvMgRdhkGJQIavc6QBgV06CD4pRzJVyUPrSS
4Ngv9SQ8EKcw1z/NJzR04OUCb6NBbC1qkXQLU81fYajxOAi7gqGq2ynFmaGi6+jE
ACGk1RyMraHr/7HPe7RtvCneaDf3FgnbKN/YbNITp1y/pADUO1UJ8uRvKUu8rha4
cxY6lxMFPcqNRZzkHRlhAIGeRNBX5r7SkDZqdMVpnY6uSO84Oo5esyHB1mvkGShP
3n836iJ28eJ3AFJnAtUREPHsmtP+qqgCXscozZ7WpedmF9rUCSxbD/vm3s/8DXco
bnKwuil8BX4qBlJYSJtfDET/hnFFLfP1ozwoaPhw8flYITSN/HSLHqgWjoG1/G5M
EvsEfFVB05dtK+VCN6L3N+zmvuUsL3bgFOq5aDZdAlvGkqVM+91X1KSpMaCX4OKQ
Fm/lX55I/lwuJTx7WRL7Ct4jkSEvc8ACEySrloZsY0lbQH5j58wz8d1LiSaOe++S
KcXLCEAbiXZDMn7Tf1dfTeFlFiGWPMv2nEk3+ypHlqsp3ZB79BrzusGnP75THtaK
JvK2kq9D4S1uZvKnOXeP/uXoE8AvVvWHXagpeFUO7dq/WnbFNkmz4yPXeeEVZPvo
Y9tmPXzDASx9vzSGwwaihNla5Rh2IrvtSZUxE6jSi05zsYLCQMoF2DDx0ne+1iZx
nOShieDVp8kIp3SXCFXj3/urCK8asnPAZxLvOHOcIIB2eNf6yUhTvo775CCPLPJV
0zNcX+2E/Bmr1y8mAPfuDoFOlgS5f0ukS4+TXT75U2Mryji2vk2BDbV/F7hVXuyt
0zFUa712vjGpzSKNi0Eic8h3rfgG/gspg4QyqquE+YAT6oXxPrjqOGxmUDCCVtBA
OJSyQM4kv1b9NE+e6dXuFKaQOMLTMjhHwFUwTe+cBxgd2eyfOt/wUvyqugi+xC7L
8hpWQ+dZpw0DjVXtoN/oFDJHhvJkZRbfgSbDjOg70YbRw1qRRDZdlqNvAn4NyfC7
v2Cj7PvC9p4HBLno2SqXZufyTkOljw1+07zZrHjaqr+DUO25wRlGDIJQu7QRPEzC
RNho4T7DTBU6a4jYPa5IhgeKKeOO+GzITzGTBZRPBM9GT9coiu9ZCqy9m4NgHBBu
FY6L8l8y3IMgsG1vv59PAKtpUAqvT61QXILvLFYzEgt/EA/fCrOSD58uhGkiXTyf
7rJujj8wOgneOd/Yjloj9tkOTrygI/qWDHoQ7O53sGqrhFo4qO196So9urF94r+j
5NbkKudxpcvutkonr3suv1RMaO85GtAkZjo6TfSPzooYGv75ABDoNG5M3IXXtu8Y
1BWroEAuWn2+1SpBPTHgEdX4T7I5JImV3VzY3h4igfwLLaPoJoTYCT16QYjDFyF9
y5AFhR4JWvhaUKSuqGo4p6x6ZoW1V0zmWLVif85vOV4DVRvjHpwU7kshlSvWP1ye
+nZ8p1ZoMEsNUsTEbZ16b7mLHX1bBKut+LbeBS2jzGiibPrvNN55RZXiuwbCGWkg
mEfsBKHXo4jSeu/5YLNzg/TQpjvM6Daucv94jcQG4Vm4CKjF60DovEjVjDKB1XHy
R4TTEdihTsjFZMMnlrS9wD9P3za75Nj012hUm8vuwgLev1u5SuAJoPchggUKdBXr
tmB9hupSyIEoEltWpX7HgzwNJXpbOXHCpTUMd64V7xIdTsXnPS0LbDffs8PSzmA1
Rcfy7QImQs+mivCVj4hy4DGQq5EKt4CddagNeSE3uG6efO2i09VZE3vd4Y68EdFl
E/m94kCCOa9SySEdb+wgX95/pNfRir7PseIFTVpMO6UvtXIwgP5eilD1m7yA+nYa
Fo+z9LV4mz367+BuNJYzXzGcucyOQXwuZMx0OpMW82daLauawxaZeSNrX8ElCBUu
IKgtKr8FHn4XItj+qD4+gw7pOg2sg5B8UQiH/j/OSaZlPz5L7CsR00CqLLWKBYc6
klfONy2DYHsiCCoKDLx7staEfpnwmGDVqv948lH7X76RiQ6+xW5DwPnFPBmTvGFR
5OrB8T/YGxrmdqZc3rEr/GY+nliBnfuEQb3GFl+yIFWaPIZjCBEKXICDHXNGGm9N
kqFN4Sw/QHzHxShKCfI7hlZm4l612awU0/jO4ijC4HOrKi1ZM84wHIIm5T/cSe4r
je1Dwamk6LbIQgquBgDLbFEtWin9darfsOlSKAKK6UFMRPp0gNZ+byhrq8hwPqyE
wwO3dzuGx5vrmQ6yxhdTvqbg9I3S2AulHyTNM5snhip69ZtbJKFePxC+XtHNBFjh
LrTl8gJKdFl1RqMdfztm1plQALYjrdHsZCmRZbi8pIG3mE9+66ic6k7F/6nbA9sQ
0Y84UmeRqVLiknhUbN+c6EHuxHxA4gbStjmIgR6rYZ2/O9vhWJS4sFmE29l9zCsk
qCGSEc3CfozUqM/eq05sTiHMgy3/1PSDORXDeoWdsWEnEcAyLtjQcC4d5rV3Yfbn
AFcqzvCYq8BndqwPzV5Mnr9AQOOX5CeM2+2KvmrR/KKF7Z1vIbdn1k/cW5+vk4eO
oLeA87zueDrs4afU6KlNR2rC9ZZ0iTyJXtN+VvMSFVY/fw1CgEp9oW1uuk0lANdX
rqaehG2tgTdgdzTMkaE+/f22vKyUAawiUM3PM/VbIqoyfqUiTKlR8fK7QLyYqj9o
jrU+8q9+dP+1efSGA/x4Vd0a8E9QYrlRhQBQZd8/BeqBr1DIuSXvwAUZCLF+/Au+
fTCDHxfZ/93/Of1yzHdDOQn15GhtVtDeCtbaHz6b5mCwwHJT5yxy2b4ZiZk49J1j
u+p3TWK3B4h6PDPdos+aFR38sJVA3+4TuCMwQXdrBDGBZ6SpdZn/dkZBBAGWa/qX
DUloQwgCt5UcoOQaAE3JBWz8LffFsNeo0QZx0hrtBmSJ9F8CcFLtc1wTLKr7/Klk
2nsy3zI/LEFu3BA7Jk+Wr3C5Iy/0kzLdtbl9KT46/VT2+HYl2fYLaVMNgyl0ual3
QDxJ42regbvg9i89cpZ3yRSM+tNKR2dUL/VYqbwjJPbTgR/t5TyImk51H7tVW9hY
a322AOXR7lv+jjkq7gbFFCUSSP3wceFqrNHdOZtfYVS/fnkraGXopJVIdvHeTYve
UVYaVT9jPt5IECrp+XQiUTLWhDwoYtITXAv/nihTJqK5OoQliKN00KiInAMLm0YM
7pvKWfjKuYGa5s73GopSSEDPEYN3oGosM2oVqxIrCI4ooIrLdSEUFIVtvQryDjzl
jv4Xomq55Vav/mL+0R2/hUKAziQcrjYZ1X3LPxrGTiUVSxBDJ6f1O7QGVDqu0eyj
coCl/uquQ33iyeLuM+hv0+QdBgQeW4J7jrH/3crwL1b7Kt3E1c50UdJf0flvhnfl
YG0Kbd9h3iMd6sY5GgoVGUHT+rYeZHggt5tyrq9TqFepgTsNae2PwzX67ZLby71l
tcm3drYReW7YSyVm5yRmmh5i2E492euFKUf3nDjmh8Q0QfG5y7KokHLOi0YQFlmK
WUOdfQCjzlTApAUA7RZnubNkoiEadw++mZCjpCUL8dFvSmwCqu2vUX9LWZfVgxnP
fGo3JZfxOP2KOBbm0SWlUuz5uQkDcC+83p+9v3H+govkSzxcQQqINsEjZ+IHICRz
uns0/Aft8Fjq+HAn/QIAcEyx41sTBQSqjvYNVmEiK1UN6CdLf/GfpHz+5iSmNZAK
QMvImiZNKSHZoZz26jjACw5A19MdknCFA+0rfA0wvyDPoeBfmU7xOgmz9Bi/n5ln
qhcloDaa4dH3qPYxpDoZGklksZhP2YImX3mEQL9F5/5rYgOSdxGuZ5PtpGM3mgMZ
i5MLgkcM4J6BKHXkTCWXMoy8+zxjEDrHdvDUX8QFTm800+3YFY4UvEN/Z2uFNE1D
dXIzrx+oZiGy8qHCx8IwFBUDRwVj/hJiGBPF5uKYLyHO+FtmUmgeGblCJUFRmJjD
BcjRCM8TQ0B9FuMGTg4MYbMcjAin7Q5zcq+53PQvJzM6Ejd7UwLG+DONcddMKrQu
f9SQtKq6csxGtEIRpByKDV1TJ1zEeK1f2tP1To7Nge3Zg7X9VKnvpuR69Dka9o/d
CxN/2u03O64teEmZCE9VSDUJnEzmahQ9KhlnsR1ftG8IXtkkS12KCrGQI+Css5AD
g4ttPfYvv4wx49eV8bVc67OgohS/RsAfxmNIrm8celWnhia/kR0dyE5B6m53lpQx
HAJ6kssT3Khb6stYa2iFL2F5uubpk3xTziN6UTnE7fn8IHhKBmn51uCs+m3l22jS
7DPOhixK0C10KvTjAmdtgRAdchclwhrmDkNFq2/AFOJryZl0R0L4indUWfb6jJde
ivSHw7voALI8VfO2wqMWl0Ic6nbZLYtB7elQJp5wszjUa2rJoNE7wG/h2UNk8p4y
FS/mlDO9Bf7YY3nRjsZwTyW+hHlWgxw/FjGYPX3R3QGD9Nlca97cX56OhS8z1Ja7
WTEuOgCcD82bftwG5Xq7G8rh8wDTvZkIMuseGgGwCl1/KNL/ZgPg7vW2r5Wc8Fpf
CvvfChp9AVS4MbqgeDahdQDxWIsvQwxnB0c1QPAlIoBqiozyVt6/VUP4cMeuXlTX
CsuM9TQNGXZMnwLxz7OXAbxOFlQf1AOSEunSUeGuQN9GL3zOAObvMkNu0hlpbBNv
A7PozJxX8grGrlJk9P+l286VdUZrYvTP7n0n6G3KeuOWOTUERlCxX7uY/0jZepZf
0gWoAA3iYMrTB0MGkSfc6/8xMNXY8hxEVElBR7SzvFZ79Vqy9yn0u2J6C/mGO+nF
9FnTXMkjhnYPhxLomuidCOzN28cXXcYTNdNgDlj8feiDDxzwXxA08A7dJXLnIOa/
ub+SrtwMzHcArRcQs45jWrjSD5yj85kzN7Hdh6wUSi4DqsZ89GKn95z9XAd7BXKB
NNjKaCRjksO6WkKs1oESNXT0LjIzOJnLW4rzb/GgHpVWNQds5CvGXRILAbhpHHW4
5P+ICmEK+SZ7Rz3fs2lP5u6NK3sf99jxeTV6mZpWcF6uyjbLuLoqR1z1W8rSjfUU
43klsloWrX1ikOhUqjsq6Pa0Y4GM3J8wjdFLTEu4FnYJj96Pc5ZY6WpENsI2xu/B
Nqi6exTBP2soZoUUHLPjlo5zxJA0j6z/0GMsRuDbMJ+mnspXYqMzvQXYiAhoKmwx
5G2pct0tXPDarsayL0m6lrwMXLWzbS8JzysdM9Hm5ESiCunFOnDJf5LNGYHmFPa0
Z9cfRLY+4pgvTOgRDWcqXIMr06ilHJp/fwYUXsqbpmpcbpPu2epvfo6wckZmdtUe
cRCKVuecnXWBE1qbDJqRmgVThLOS+a/cG1AzS1HP+LAlUl2QQVl8C6UTT3MK4SVT
tz4CGeSrSNl4WV+8JVBq+gGIIZF/z+T3BAYVG1ZGOFnvu5BU11aOrK8nWXEjWr3/
O0OMXzcUDSCqlI6xKb2OkRAC86GpqqziKv7WkRWlVn4iWJfY0AeItEOJBsuo85nw
URIgNwJBovqybY0Ela7U+umlKzAmv2EZ7DTN8ClozV1AsnUxeghJfMpbvEvh/gIQ
TRb8UVMseEQ+OffTbx6JErjJ5+jSz64LXrzcYvOH8Ji+m2yPkswZncyhmz6sUMAJ
hLNhrj5iu7bJc2KfvJOgPX7VMi6aJ8S5y8rgg9Xc7E2IGkAdmJhm/xxlYRVKkeiq
FkekWKGDA1XL2RHt67uWEnqhmTNyo9b+ACLkKDKRq/RbBxsGTFuOlcm9iOiKBvvJ
lwnka3nwYZ+ZlZFakSIuC9QDOXDogrlKlrfxZ2mKes+uw0P/3T/yqjTLnrJcvsuS
GknCKlY1JiI5vJ7cY5WJlcau7dAsAbWpQBtrZbMZFjuMbnJwG/+25zseYMl93yXT
Q8ZLJepZ18rkw3DTL99ucRMMUS4UOwAx3ETx9BbLJ6HT3GvOZprUn9UvdsBzbw8j
1eYL7IMw1s+vGaWfle2UvMI0qV8Vs99UH5Bv2I4/3L2JPTG2T9+j10bxZPP2dIn8
u8aF7DO3kbugCNgX0eNzmXdRpZuRClTPQntvozupWUWRVg9KCE59SKO57z2Dd4wr
xarM598tNlCfJt/ICE0SRM3ACvPtHHhUDMkoBP2EeSxfotKHXx6WslSzUxll9+FC
1sd3CsKqYOj8IeMP5G/RLqq5e9vsRydKP/eljdO7qLmieeHTeXa4I9aG9z24Zxo3
PPSktlimbdfgbAKlrpk2LFken/qm8qclGGEvUQTBCut0gZKtrHU8crGo5nfwglYl
SyXfrc0HIBY/sbcR7vqHEYlt05qXKaPCpDIxh+gbO969ee/0WG83WYi/XJVRXduI
TcxsIpd5US4a31ohvyevbVMna250GbbTYOO8gzr8GOy4BeoCfhuz76UDI2sDB9mx
/2BXm/uZrl/0QQ/+lCV19HFHDDxNSphshjnnyWS3qKkSmmIK166O3NfEhH4OGPha
zdYVnSj1ISYVpGcPgC43VKSDJJjyaRQ03eg+zSb5cftBPLtYHJKo0rNaGy1XFRcd
7ovnhHxUhloWy7CAVTg6B0wNtB/3ITPNu0OzVEhMDxYKskccnnK9znbYrZNUsrC3
Hpnr2n2GGqDok3futYxKuNyyMUn2UF9SKPOccvjRMgfCPFGkjqHbCOBxXl90gEpB
/GZJ/lLFIdr6HgmdwsKngsaBPK3JPz+6bscApavXmUnMJr1Nwhl/QD/3xC5wMYb1
XEYN7K7PSEEXAFGCO9RRiP5ODAJyQemeBU6ge3wDQcpucIqWIwx4dByVY9JUUovK
IrKtd95018adRVYfckGxcNwgZ9iYK6IlVuM9URnSilnSlWLdexLSSePSqPgruNQD
RFbNcbc+/9TosexJpQMX+GYwRkAsHLKF8+LA2M7NThphjHM2YlC8bhtbzaxFoZD8
WEwy4ZZLiCYZxRVHrjtJoWFjnPHtS46BWOJg+PG5fQfO9COHep97W4CByCkPvVrP
6hJhtGp+29fiuAklpDQrF1AvRW7lb6WoN/GjSKKq1jsdssQay0vbRqqdFCFvw+S+
F/0AspHvSbCIAI4lUBK6Z9yIheM0BL5PsL+p2qU/TKxUv6jGw2sUesVzEXn/L6Bx
UeRX4m359lZC+CPBvWz5q1Ful6t7yNoMYrUY7PMDcHhwCO/fYt0MZafKl+QOUv4T
lZYXxaBhqr8xU5mZpnBXwRNMePjmod7ZjlGKUqyJ0wwhHbpPJshKLBnga4kDLbtr
1ICpLrGMBGgYAjNk3eegCN1jJlNmVbfTbls6LoEP8uxDjNqH5d/wHiXgKgPXg0lI
cJastNKS6n4IHj2KhECGgqHaNp2a/GYQoG9DFzHo6XI1eXgXmA/QvfXaLBCp/P1v
i5PyJCYEjiOZN1MWkXoV5Ew4i3L/wusJyEoAhgW6gGggv8y7/AX004b6UmnoVMhe
nJ+yJ8/Ke9wR0mr/CjqzQ8p5J0KP6Zso3Owi/X6PGiadYIBORjdk0Vt/WWSerDvR
Cq7GeBVXg+FZyBlG1U5Wol7ulzhSF1sXEWT+FWPtC1cyk7xfGFgw2/TaOp/CPywY
fmrSIzw/LNk+OFypThOAWXcvSrDhpEPyBwU7yuye8ru3ZDTZJR7czgEacjNWx1+d
pR7lDTbxeZuYnOhZAtobFYoRt7Yftc67t0xMeReeWAvBj6ac0cAVd9RA1UVok8Ls
zPiEcgg1bq2AfFgQdkHrMGszBM6V/+UDshSBUi3V+in9nY+2qeA310aT+4Jfug9d
8QuVYybJNtX78Xka0BW8+wO/FVYeNL0b+3ClMOS7obZiToamR8PGPKOK1WZs+m3L
Pkc8eIciQM6sqNJPHbXCSLYouyeJuOjlzDDZjl25zdmmJl938ZrPADVjvRUTnyBW
kh5kAenvjaUsbRkIuXVTURdVOkpFMP7x2hDfl7rtTP1OLwuAkEflxGBvBrW+QrMh
sFE33QzVZg8+90dlDcvlxbRiAMewWgJO7+/lQrjqzOEB4Bj75ekSZqnO5cbkTrmj
t/6UE/VGAfgCWGIKNc0X2HWRg1aiR1xiTbI/vCJYWSIT8a85bMqs7ZeEcQeMjL8O
OtqhbEuBDNbch2yKdHAIg6d0oVxQEIIbxdZVoPCJpCLvkOPPBP89parWOhqcs3uD
HjQCpXHaaTMoQZPMG+0QjcnHqEVLmwW2J1V3C5kjHDRT/fjRroXOpKgReNCBOzvD
/0rNwvKVA0/GFJWkj2z6rGtmRijQiAkSSQun7KWxUYftW6aENXk71mvJy5XUxV2k
qxiiZGvXQ+ZHKCfuN9SG6uRcfkDiHcyvWoEqPS2QrGPahiTYpEzxLebZhwVmfbdY
IE2frhg9Hyv60bsl/XIdZTZmgxlb1eR1wGaBEsgW9nXNdD1tf+qUVj2p7ZuxnwDU
aqvwoLckxXHPUtVfrLGr86Z1KNAQSYdKVoIZkHfxgPO6VzFdXPXDgF+pE+P2VmZJ
RxAnNZh7/9NFKu1yJZQFsZcAZ5hanbchuQ+nMZWTrkwdY1CKQSYFhZsxekuJn+/r
bIlt8QyO5GdcmsNxptEXRAF+RARZ3Ku4EKjiibdbrRXsx33uS7gjQRZYvPAZKH3e
NTmweFUrPl3XcQsoXgQGnfHcYhaoST4dyjKXpZ2Bc2H3ysqLiRdC8EnzmSYPndBT
OQoBOBPWZ8YrhW5FLJA6/d2YvCreFXkkfuoqBXESoa1Fm6p16BJ+QHXvEAkKsbzB
bpQGmYbS9NZgss7/RWRgnwHjBoc2tww3ruxvXjpIOR/evYqsX/gURr9hk76EaqyJ
bRsyQl6BVugm+M3uY22nZH59VpKSteVRHAx30hAbUx4S1xlNTUGXHyibsONoR0+f
Ak5kIMQU4SUeg/lEabuRBo1w+LGSWQ6QDnW48DinyfECwjeUvKRlAbOI7Bza8TUA
j5m9FADYXpdInZSlr4aIdgJZZNBMrF0+D8w00sxkTND6JD+BmUQ0Tc4ITQLTREfA
8TtrWr5NcVljLVNg3PMf9XRpRjVBUvJY7Msoht47slkVbYs7dJig2AqyHkYWMwBr
e12rU31ue0MEA/hCI4ZHh1X/4igU+8rKhUd5NdrRt4GKhoHRBtvt7pdaxvvxbwit
GLOPwFQzfTbeJCyn4VHI8hPcc/AtNsRD0unxYuqX4cr142rjf2DNev7hvOPn5JBf
SpqaeoBJUlmFZghu8GPJp71ChRXGduZb2qJCB2fEqB7T7uzFpv9Nsj9TcrZpgwxg
rPv29aMlOUvqPvp2ocK8NfZcpSdwyVMHbnisX9wfQaA5WHATIzsMS5IJIGn2RHNm
rQ6R7CRNdyhkH4W9YYj8CN4SSSlL/eIEhmNAKLZg/7ChnetfeIFK3q23iAb/EO5Y
p7GAEt3wZjkjXZUmhXP0ReVJkdCPiqscHwDpYGvckiOeGAv3Q+4ysoVaP8eqQFNG
IpkyEQCYzqn3I9XFhkPLjpD+p3naCA5UcKPvoyKvfN50VA4aBKsDILx8YyHi6yU5
LA3OeeYexMvb/gDWGPLpeEWF4WcD5rU6g4SpPSvQKmIxE26wTHFrQ7VUo+slqW3w
gsLjG0DfX1uCIA0eL5hVudezo4pCseWobapJ9uK8uSMx66LKohJmek/tmNDbKQGW
7CHSnfnjc4R39utF3juhsaBY7nf7TVIuq+9IIPvSvPT/+ZKxCy37CqrEjlKPOTTn
d8Jc2NDOzXjhCT2edVdnfLvLekuAYcNPHwG9jWJy6f1g7teU2GG/aZ/9kN3f0FjR
30k2mfq6oP644O/fJYF5hzfnd5X0XjlGaL+60UYPGJKMAUfL+z/raOfadS3DYL4p
4MsthQL2pmwhsqC4lHlC95KuDamjGgYn9WG1Fat9Ez56kT4jpebeKvQNj7S4ncM8
4z0mgoChiB0XojKEvwcxHIYqwzS2WCgJgevn3cUpGAEQ4VAZnH6eQ13gDfn2DdWZ
XhvWBsnhIlGY3OzhNjCOrH1kKdCL81vGxVe0JO9EB0RcPP2E1jWxLs6zxi2poi93
Om8L7UHknMCpuO5QrkbXTBeMUrGiqYdAzVyB7qDidF0llmFM7Hexm3ZO941gm3x0
cjnS13RxKEZwiTvDXTMaf4IuHnlzpDTfKRAurQcmS0a1+Az7dH3MPufJKUduApjh
RMo70rpbEupQSNiibvJNA4E7Wckxra143S3gGVUFBRrpF/dxkjoXGvgKzH68A9oo
o4A+TAvJH8QT4VfNVzSXcStmKbelEtXfeiE+1Bv6V7ZaLsuMjpalGNOTvVsxIBRN
l/WtXfltOGhW8PVFirv3vjjZ7vcbZ9lGfuPktSoW+wFLCGMiSWtsaZIqkAe/Jjg+
KF0QK0nP/Fb8DjcFU90yR3hYfwp9NZdYGtDZHiqZNZ52hs13AIIDQjiI0XyRQFFy
JP54GNQXonD+QnoHhgzwOkoIqJ/PQ0Xdeq9BNUolPO1Qx2EbcGr2GJxN39xFctqz
G7GyvRmaHoE5JVa2+TxaapYMs4pHwENGNpm7ziSHEmBOgXYWCFk1Gvx2KcmjEJl6
2y7i3sLYxulIE/e/eVa+ixtxSg4tjTUXM+DZb+hkTU317NZTjNP63iLcqOwBdo+9
mGfBlgfp82OUuqU69jZPZTo0RHLclJrVFpUUr5c/1d9jKGHYv+U6Jxkr1o7aCEuD
WUC1rakBhVyEx8SDfd6NOIlH1OshZnvGFqFsxf9N4KWzrFodW0DpQoww9lc7NQWR
TBDsLbcrPGLZJaxcw+oWdWBCSzdlThR7oLCRWzwHwHbiYJl0ewylcRnaxnCDTH7l
O6gx1xID9eQPOnTu7wLAdJkixM71LqvWiLI2MFQOoDZwBx4rEeLrJzPOtDRfI8Zi
0bbdPpOv15Odg85X/0Y390lQPINA4PMjaNnjOe4/oZ3RTRqXzHAZ4t+oXq9RNvCk
zdy7neIlkYs2d1BiBFAeAloooCbLQyfaJySrEFyp7nywoQZwA+/tWYfiBMmVIAqN
PbWrIdnFSeps6PrweNBBwSK7Zq47p0naQC9xP370Xjuij/9sqlweiGq3BJsec8mL
ylJeZJXdC/sXAvh5Smx8BY8qEwl8g2n8dIpw4YbJ8F9lpVuyqh14jiw9kSj5Z9bh
d81kN0RgK1tgZkpq1oMZHRWyKG6aMaAAS3sYyKNJ/yayWgxQvePurBIhcpZnPFMW
8tcVW2iFkIM0bhDjZNgNn/iky+dFRaWDxv2XO0S4I23sFCihRpy/ZklVv4/FGrJ2
4fcFAV8IpXShPZsy3DAviTM2j4OcCvVyFe3UXh0YQppZrMw6CcCmSY0HKCpo+n5K
4ZB5QBmx4Bj+4nsqtEiMVAVeGdnbODjS6BLiT2UpD4426RuYk3qHcSdujq7by+ot
mo9k/9tZbhQEgUuWpqXuTGESo/2nPNiDDsJJMqG7Um8GVEpYx2yjH8UDBXgtWQf4
goMufOwMZmXJw6TTQKxVV3aqEYzpiNkE1DkVjF2wPGtpOxvbHvyp+2e78cOl9zm7
fAowHSDijGupSU9UQniSqL1pBj0eD2bXgz0gidPnkP6SlioiDSR0vaSfdrei2BAd
pRxRD+gvoFSPBzraVUHg6VgVyPHSptLzepgTNMfLhV4Ki8hfrv58EoyKvjtXXNc2
ZWB6PRrb6s/UVWCrRalClRC/3e1vAq8tB0U0YzgZaJbIKyK2QWU+7wTpPL31a5bP
rjyo07YwOUP+xhG8Fc8LSdZgRctKpfA7+eTVtgRbYPD1eopIrv5MNmoLSzA2Q4mD
jDlYiFvQDHzFLitRkoYyDv1b6xo/VQgGCHnbt9L62zXUhdo6FS+BzZA4R5ISoc0A
uANtE9Ctd0Kv89sZ9CK2ug1Un8DhH8L1pFR4sX4XeNJWBQj9sB+XtHI60GK8ASAH
exukBBARdz/AiZ63indhzFr2GRFDpy60S3hdvRNmiSQxo+6XBbD5DWMpALRRdgrG
iftNGDdqH0h0dDleFNeWVT5HDYmX365nZokRoM0HLcrz4UDLyBP4VxUE3K9fpypg
S/3l5SQWN5GXpCS5iUzuQBpirjYzUSkhJNmzfGdtSlHTezJZ+IZQy1v5OyVxSKgI
tyLBsM3jHw590qCDgmLqiJ1srlL/yhLa9LlvlkbrN4yco+KTTDzmWHUsFUnrY9RS
BkG0pt8ryIWkQfKb34bfDq6iEzoEOZ+NgEqwnMM4RMO8N86toRilWgnIWQnN9Dxx
5i3shlQpYyVM3wKfV4OIc2rkb9u03WFs60sv+zA37Mt76u4dBD5p/T54hdcXy/XF
HCKWJteI2IFWKflKxC4R5g6AoiuRNzuDpRB2I4FahA0waiOXUmXbexBj2ykpo55c
kOF9GZ8WIWnT8GctQ6qbiGeQzLElSTlCziYOcirZrWhBmO0l8cbVbQFasRr3gTcF
ekuK9zbwTA1TuUBXj7aflCP9w26QpHCJZxPLnOFeAxzx/fD1GHdYk7Fob3kPIO4H
qhXJO3kfpVvp4Vz8Q/SJdaIi9HuqxMJCcgVg5bKL8B5qnR9ySFEoYTV0jGt24Lh/
e/FroAf2i6lkIRxwarIkkXbzt/SiAs1MrTiRIE3YCkccyxeLaZtPVo5bH3VHp4qM
hwvYXGngUZ5pcSaNf+ivlvnxHunqBsv1IPDV8oIRhr2mfvQmcQeU1CZdxbm5PYPE
xwQzz2BtJ4BU7058MHApjUnOs54N5zMtXfqaGnQVHC+/FS0/jc2eVkr4dk/Ikab3
omcEc5Q+NdrQgpVTLAt4gzIEnLvVdpKkC1J3qaPMwgzOTvhyVaWlfnC2d5N320H9
RPd31wuJXqEL9ohxK8+5C+AFWTAszaLI5nYc5DxDWdbNB5gjSXP3M5KWcLGEHz+h
4tK3Mk+d+GGw3f4NC5seDJkfXjoc4dkwq5wTlBzwTHLN9CIJmf4PlAKzurjuB2ML
fQQg1oe84cO9LgFfABsXe2GR42WXXOjVfJQUG8kHFeP3P0XBZqkAebOIqc7TZkVR
gC+AJ3a5aU2+0SyvGxPg1AP69qIoieVgxrxjXlxt4LxNXhsPX/oWSZf7snd0Ht21
Rar/jupdMYTy8mTiRt5CtmFQ/5MurH/Svqcipcb5Nbuu+kchtaKd8ifnU7UrEYUP
kpmmuIQZ5Ed+x7Vzjj2xwYnLSXLS18xdNTvk18USmvLgxz03lq/OWLBuFMPOBTC1
vz/UWfRemCRn7JLbAuJn9Res86qapbhU3frswOakXl431kZS3dmSAPA4DWhsTZR4
kLPtuDoA3bqKZPew256rHAyLtm5jklMFjO1m99tFOonc3GCeT3qdbdFVUAzsXzse
LjzZTyplmSmNZ5Jsp2lFgxCLKHKZiZ3GY8eNSnKRMWryoBlci1E2UPVmE4DWP7zM
7TR+F8wK0o8WesmBteiFVyTtObreyEUlFBBHuVrg/TlH/uIUr0S8PcSI5yj0FfyS
moH9V19fYvXUfwU6/gHUZRCSQs5IvlWkCDlQnq2VFnfQdvmhxAxhfmeCXNpE3mm5
+40xLFk1hR/WG0zkDuqsZctOkyMP8EwOMWmlbsoJ7D1oTe3Zoswz2FL2lbLUZF5i
iRF5kjDv2IJWyq7ZQbtga+S22QHiG0CsRZu0FS2QcIpL63vF/g/Hg5qlGt3JWDWo
88vERKqU8lOMKGVnkhyLZW01520WDyjXs6UO1Z9fMSgVmJdBLxokVSfUX04EOvjq
OJFrcwE69YGC+S5Up3ykqbitEFsWj1RkKR7OABB8ORqHn3Zl9CrTPp4DKF5g4VlP
+//10AGLPzovzB3m/DoPVLSZtalkJE7H+Zi6UIPO36UmqmIEPJ2lNwhZtL2OCtDo
lesC4JmKnUxTGPQeryZCujt90+YgKL+3mzb6GZArs9LAaGhDDx9pFCvoz7DP1FYn
bRCOZYfio0QMYC2H3bn+QrXKRUrT0emOjtAguxIW5w984Uy39Z2z6kQa5mMEszoC
ecA46OZ9vFTouEUkz5QbxTpopsVBPQwKL3g5pYXGRmR8ODuHJoaCQqkBALiEjVES
u14LOGUoaUxyCY0S/Jp/tHLNSk29a6fZyMsK/73l3Ba5n6SV7thfXvNt1qJe1M1O
ndh/Xvheiou9gidROvZ4SDq8CY34LGTL0UIbP5tfoGbe2X1uM2nTWWukXeHKRBVa
jr2kh8gAWZeU5eMhVEoqNtiQsRozzekGh1dUVge6J6QzNIYu8QtVHoLwVVR6qVmW
F9R6qKtwnBmVUgPgu2oixpoMWFps9vRPxMWG5Q2aK9g+JMocP9vENurTfKZxXxPi
wFBZ/pQyhgjilLH1X9vB5FOWAhmGtaI5GyzyI6R1ebNuUQXudT7m8HEXlQLkd6oI
LcaqWQmpZNHvb4PAUNzSAq7PAz0Vx8mFsmrRhcnd1qICZcTQb+K0YFzcqmAftns0
3S8uffQ5yS/wVdnpPqmfvh7tFV08ub1290/pkoa4bSU4rn8sseGunORKWnIlLqEN
t3eIJwyuxjUadB5EAPDHaXGem75PJaa0T8W4REU9vnPTHJ/Qgpx8lMQ3pMat5ZsY
fsv3P7refzeOOw5EGparz9ZnAuevrMQzEAsOpJLeT8+HFEJ72O2OOfoa2ds1qNq5
6rLxu29J5YDuVC2KIgSudzHmoFAFrTsqF/jZ7ZPzKXaRB18DsE/zyfsA/vol7yRU
Dgh5IjZ/hRaHIDYv/hCXVHhma3l+AEVvC46HC1JsbVhSwRB4oqrHkVYcFJdPYjo4
DfJFekD5/LsjViYkIuPekEmO6QphEwXC+QDVAAI5ggmN6Dw4xx1dMXRu0LEky5OY
UOM9KG8xRZCtK7eb4Ad+C41zORLwQu9Y/FFifWAD92dXePHZUSuz2WmITfnOeoTn
Eyoi7MDpqYKoJZpS9x43oR9MXO8tV2MMYE0RHsbUInWIgZe69K8u4yODCZwdpha3
lM6mQZ2MrhSMIKHvTFJN8gW3hkxe5tovnRNLMeekZaOrsaPD8SaOBSmUd6yIlBk8
wF/eClparA/HiFXf8VlU5Ohxf22cpCGbHgIQ9fXvncow55gCysA815PUGr/8iMMA
DvzfkOUCzJ/a+OTtfuQHWF0+2/zEo/A10s05qirlI+XY3ojW6p3r9mbdKoYGi3k4
++voY/eLZ+OTVZ0Bz7IacUZKSVr8rr4jPzYhqq9XyZCIOzF2glxtkLhjj4SmN8T2
En7I6YuNP9PwEVKOcrZc1ce2boYhHyaHC6xgKDIXW/2yVAiz1FagxBOIDAY0+96S
sWk95kDVJj1BrYSYYNgiYClcGV35x3NqrG5xbB9BTE3+szqSCNTBqlDAdJlwD2uq
w0e0U7evkWRMXX7CuirfbtGBw3+5Hg0+mxSohBo1pqqYSdkxFj6O0xgPQgNPS23d
ZtF2WzHs3Bmlm3gPFECT/fSEsjbjrs0C3EOeCMrvxWuRwJOav3shmT0BenTdSIUl
T+1/EQfp1AEXEdGA20hgk+YBPk0A+bFh+52MUXLaCODNPR78HYKOVxLdSXK1wfAs
/CTcfKXLr4YsDSQcvCkFBwwC7ra2a8gyx3y/+B/OnRXmn6w4MycN8zuD8D2U0/oI
fm4EBlLneVCCLi5qgCyNAzbaAy9IhCvUMzDgn2FR27s8mUu2zvkNA4bpv99Cedi0
FfImxAVP+qrCBSbvuusWsRX9kZDqSggQfdS0QKuoJEZsXIYD4kSAcCT59IhS/w3n
Wlwc4D7hy5mJN8YE+NIqg2duYVpue9Tmy+nvpyx9zh2D8r6kW0F1jZEWp6vpp7OL
E7cc9iVuBKospKr/mxDha35HnjjJD39bYl3/yPyQodvcYpIHnbBYV6e7Qv95Hd5a
NevWIEdlQvfvEstvVa8E9t6Ym/lEY9xDEto0u5lRZY9CssAeVstX+fbfMxo2L/iF
iMf/oJSQp1hTIJDbV/AMZBR+r0Y6CZ9X/2TLw7/mEzVwS2SVlhKTwS7wNde+wysu
+Zx+REZYVyWrFr+b9/eniTUYN/KsI5Pzu0q8kE3TzkwkNd9rTW53lfj1g7kOaiv/
NrNCwTq/6+cx/YY/5N+BTQHWdpoX6ZxUgeHZeCJSFJ/A5dZ4qagZb0cNZFUXpRl1
GL1OPslW07SzJhRLF3JK7XFlGfLJxuhi+4HuhWsXNFCBwVcZOyvgdgIMLmlTUJUk
wWqXhT6VdUs2Pg51OUU7OFqGVmKXkvu0pJA3m9MUXfXuB9CBUrdU+u+tw//Vyx/T
05A4zzy9gzSi/IscQ0b2M2INMsM8jfvM1HwyASCQYhckpgAQ8xoivDsM+lCnJHCO
HfmY7U6T+TA/eBYNnBUh/61QcM73IyGTbvkerA34zxIrdTKEH6e6U1xgzJMywVu1
U3tyF2PBftiEER6R1VCm6VvXeC0DfNpo44PrRdvP3yz3RYgKAdU9E5r/bPHT5lFD
qOwYEAryF3grSpABipWCmuhPRku8MZicBgLmCn6LXfWeeHqShHaD/d7MqNhrsu7W
XMqWlqQGrCqswa4M4qRqjWx3b4r1j+a7SduiHgDFnU/wIh4NWtQCaSqgX9tif3pO
6piYUdY1Pd7bsM7oWxohhFZtY1sFnlCQAWiR8fG+eiuWPxDwsqtXZR6vlelnWfJK
nQ4Gxwtytu+wAG0y/yi1DTPW080Z/ce9IYsj0gYSjp4SeM7v0EiHp6esrcI2Wchs
5e+Qrbo7zsQ24R3a3x17YgMzhJHbVKVDY81wf7XypFuFykgJD+QN9IEb8Btlv6Lm
Xj4rmkktbk3NOf+sA+PhCYrt+L9YbbaAnDc0DDu13T7NPGNPVWaQ2KeJ9AV5Tpnt
3Rs+k478U6adF3dneMy3M1UZzRqDmwaeYgdDnGKXkZMGXwB3/IvUqmn1S/w4S8ra
9Hv/FtngblqNAtoJesU8jT60dff6CEf8HMiD646vPPJvyvEcnWyA2rRam6emA3Pp
xtjDzR2jI+L13WblC0WfbCQA6DquI+L+noiKLzVCaaXWz25sbhLEPNFAxI0Dg9N4
zJS1lzGn1UDPrh/b6JMuLre9jS4BIk50b4AdrT3WvPabB5mHRkuNf3H0JIXm1K0B
GizFXdoVfIFAdsf4PBvRBLOBmFCqX1ywRnuK/GifZptJVzV06UIFYBPs/sRNZTZa
6I63ipY6UxH+Whf5hZARSqpcUmSlIAWos+jQfpuckacuMmo4EAySexx8o2cnjlc+
K/qxpHn+/3ptKuh85dGFHL0DnTci7V+kjNr44RMsIWorEclT1DQbQ47bED6D8Hew
oqr3FNmFpdHS83zC3QjKXACQ8TC5CbjishoN1Y2qbRttAVef0XDuYzrFKDEatebO
3YBU0Qp7T4kH73gLqJH2+rGbpFvKRFfGvlvRvR0PH8JQc3GTEesqJU9b3VWqb0NN
wBCaAy9pTIlsubyfo/laPRjMFCeJeIT4tOGLZ9/p/aY4mWxKYjsdxrAGkOQrn9Rv
hEuJ0BfySeztVVjkoVz8aNBYUFseiy45UBNRHUwu1pWHEP+fiAKzNQ/8f8XJMmG5
7A79j+KMnEdZeTHYBkMcoRmMaLMXtLjhhKmLJGqrtVhGRvXo+uQ0dSE5jKfN2yHw
smfMxy/0KHN2d22jeNLfhLdMXUJnFNTeSNspF85etPiwPOij987h+oUUvWkJoA+I
snv+hCxYb6MGfHkB0GQ0Q4MrivJFR0PF89dHk1bBeYte5nLnk2idfej9+CJuwnr9
fPWyRT0fGXiqVQKsnGO4gHEqMjE6qGMpM8ba4sKFZwi9kg9IyGoOs1Lvf/idD25Q
3QygzMomwA+tv8vFS7G5zymcSFL4Y8ndg0q7p0jaPsLQTjCTGZPUIGM/GWk+eZLq
7GqYv8de3V7Zi6YLtRx7qu2obyMs8FMJOdHWW4Ll9qCiSulARGriaLkjD5EjqGMc
CayBLwlzUTh17l9Rpt07fq2CvsYGi4Fv+AKp192oE1RfS5QkEo6je88EbSl/xX8c
lvEpxykGjPemVBYKn6UsgXdiHmPT/s8VbrLVMWbkdMvqCz8ze/EJzJnHLr2+jIq8
lkVChezta1E51zAcMqyBVQqIM92uRlE4mq1mwGH8tUk7FoScjn7m5eEtBcFAOWvb
k1TaG420l9te739en6lkzPvG5vRewypnjVGBLG0wHa6qVz+AkzKFaIdP+g9axU6O
MZVgQCJzziaALqaXpiE90wvnn4b27lIFS8ZutF+jBkSg3cRg0fSU4EB9pJXGJY+2
4p18XY/TDGprlOtBXBAO10w7VzeidK7iwXV15DM5k2iPIFI+1P8Ua8Kl5xpvNpNg
BUppYXVEfH2e0SymVU9VfVLsrE69HV0pJb2P6pP+OJanMPXLSzECx5i6zo+KtsPB
ZAfhVtqhlr02eVHjDZDTvSdNxSdGRReyww2PJpscqzBUIHj1eNMh/Vc/Yov3L7hJ
BWr+tyYspdwk1pANn+yLL4gS8uA1Gbku1BL8IiBrUFJSyGM5HWV9kCkKiAEzM9+H
jdyRiNnoJo1ThET2KETb2PEiXgxPCmPsHfwC4tHnq7WE+/M0DurZrMp3gY1Y6tbG
DAK1fik6OfHRpuHe+4x3iJlgKeIu49jBce5wkXofllct4VqV4JriEM4MVhmd4uWx
N0aA79+iwr9kBfxlPkW0kF+uBuftkUOcHBt8sX39gM7NVmeN+Yz0KgeyOOoNfd/U
Ixf88KzmY1w3Uu4NGi4EO4IWrrGqGSp1TELOsMi8uv4P1A3n3w9+7kYVbCFHm/3L
XJ2SpWCh0vx9bJp3FJI4jgJ460GaBIvILI5oLdDPa/eXltfTM4KSQTk4tclb8/DT
d0l6wgvmh8b3gZD22ZRV5C+JDOoAqBL7OWiMohc8iSaBhXfJOBh1+VF6w3cE2uYk
FtvNF7miytxucCmPYxQ3IIUO8TAHAUw76h5PD30ASQZNlzRWnhJdLA1LdLLlbYHo
CHnOazhxweGamAfzZJcyL9hVlbAWaiRrKp2S+nGToOqiXTFYgb6vxkBa6MNpgJNb
rG/TIfERVJuaneZD48AkSRRH/PZAeaiXpA4MOJqfeGKCCNqLuCeqwaCZPsAxUnhO
yIrUbj7JooK4Xr5iLJ9Q1pH0Z4XNHch3bab1Ncyd4nUm7ETZZziX4VdrqjjQmzg7
2l0dyICvrXn2mE5JKKI6caRDRSb2mIR2bK4aZzoDjG8bRHztbFyRisDTJ6OSAEbu
/I5o47aWP96bKryKLUupCRcbpeeofoEGUmCUcJEeMspeUKT+RVC/reYWTTGVMCYT
oj2BjCZF4h3VGJNbqbK0IvRYNLfwVv7v2mebri1WNSn4VLL7bhjv6iOfgAggOqvj
2VblgDzfBryoA51hXp//0QUhkA5Dbif1xolvrIFpVU6ZW1OmzVOa0SM+Vwlu919O
3QwKYYqbsVhXZWNeLoOObqxXScsKEgDWpvpsOmoZC3zW6FFPHUKsIfBtwTim8la8
OmVBkjNcZlM1coUHK6YAOlhv0UhAv+6vkBGcNVOu5Sr3rnGLN+bLzQ4fp5J/dTm6
Xso4zBL3kjyR9nwOtggeSX2mBXxP37oYXmzeUP/kn7OFlhKDYmm35CB8BVu9ZxjP
4mccb5qRZUyAqI2pElKNWtMe1VpEm8EjDx+nipXXDA6i+mMCs38EePnBkytbbwH6
yAL+GuU/uBgs/3ZOdxe5M5LrqQO2DEqFWxNjME1Rnf50XTYHR8eYWLbBwbTzyNCW
OeTi/0by8Bpeb7nBEQknS0cUg1mjIsXVSOd+AFIYyyvADnDlbNcLo+Bzu7zOoVxX
ieHXuz+r5zm2zEJ2zP5olRmArxemVQ4Q6gPJKY2b9NzbsOdVT5jVqFnNhajXMNMJ
45Upq4YeeANQD7unmQkIVnpeH+aYH25yY3d82qPvlkc9RyzSMvwa6ArfDjcGwPyo
CCu+hdL4FYd2x7UmbvFCFpqhgS4JyAxkPdGNa5GpHT/5AcNIfB1RbIMDT5fbbJou
5nvDMyNHrxPznKt/zOzwbgEjS0yhk2pcnlS2qCx5jsN7S5N3C/pIvoVynlDPLv63
EPSkVTVALyrCIvw2ZP50xljyxtgayTCsq95dGenu7yLZBTsxejVc1Vwt3VVXffhu
sNUYLZUpQMDLQw4TBMO6C0/6ZqWGpcBSQw+7FXX//b+zkPIDO03eyNV83eAqa/4T
kkad8mxJhz6sNzmtfTeuNVzGmzEDRVbz5aZrNb/YcpNYY1VwwnlFveviOKsI+qmc
kcLPuQJQReyLd+kX1njoBr0sYQpyb9RomhlOAW0pnqokpWDZhFJ+UytslLDuuIm8
eBy4+xVh9i09AOLUV6dYL32bOzNNuEmJctTbFnsqSGzwa7k45SOEVzaWbxOgz9Gy
AkyL/M1eBO3Zu2f9vwMyM4NaAdMY4kOFpdtP5F87gt4ilfGM+tnWoUrSREO3g0xF
C3vx4C4tiFheA6CwalQuz+EEa2wEKbBMEnozkwfUawTcmaMR47AJXCvKjk7mnFXF
nNa0+XgAk4+tk7lQiozne/NBO9oHxS2rqUEM06VayYwSuFX0z7qxbfzck08sTrZX
9IK7mKQt0xbswGcte3jqadKkMN3zxUIqvOUNkHf9cek62izVVKe7wZJImLH1P7Bn
gFEJmGoZkkOxrE4obVe9/dXNqEaCyXwx3/5tpQQ7jBuSrx20EntWybD3w9WsRAQZ
uoHC3PXg8EA+Fexz+fFOW2n3+r7P9LXl8xTMpzsEzFdF5g+dxZR4cGmOkNPg55fV
jmZQo3K6WovTKaSr4bpNAcwXGl9Qsg0kWGiNe5XseRHbOOAbY7DQ2CiESo+2Kymy
SrlbmCGArtlQPwY/qrJuBQUgagmB9uIXfk/603z5vWqtU3ggTzplvx05nOP3KkhE
yZZqmcTaNyijSFj3PyihWjqEL3ESXpGh+6xd8HfwtZyLpmftK43J9jIR12T7EIJh
ztT5GNEXbyqwE6Mu6vSNwro8dlS4CMRnZykXMIzf/RBRrlrlvHD7fnetaOZ5ogtS
pLQj3YSfUQ0Jz4cmMSIPjpGNlBPsabHcDvDjw3d4jizfIdCUa7q9gMmh9hiM/Qty
G2aNby6nTxhbPdu4F80wbs46dKHgnpL+y3vAbbfYb5UYVD3Z2bhjg3j7XUvjgso2
GG/FmC9Eo0mu2OJ6jwOfAkDyiv2pN7pUPBsJaAsvyzFVxLLYhHbQIaXvBqxlMCxU
CZbOGpoqk+agv9+uY+KpvunDKWdTCxZSCjjjTXq+NwfsbEZrjhIFIyuJzJltLD0k
pvkEEWZoSNLfZ+YFJ7Z1JCXsy4WqBMix/pbd9SV5bjYAH5BLOQ01VNbyIwLDRFEa
i0Fwf6Nm+x499gm9P5qlfZn9qTKXMVGQHQjodA7J6rKNLYCQlQ7l+bdGvlrmnPF/
wD/6wVLkmFx+wkl7Xnq3otDrV0UckWfptav5kF1spHZYAb52+t6h4/rgfAUgQt2o
FLTx2IzwlQHnRFd18wlhqW6tH7EySdUpESsXjjTPefHVBAk31dpP4K/nG9ltgHoU
CtXZ//r53O+lLoj9tsp0m7UQcalUkQRRHJFcNNWnmf8gryk4293Psbb/IcqgCiDi
Q8Ks9WEt3OZlz+P7ncEmlLQTgpetWZB6+2U8/7OaP3RLy8nNLJUvrdJbHHRJs9fw
zVfbNFNvWUvwIP5oeptcvzxEhTHZcbD50ECOQNuhZwrBcDbIvVtinyF7O+dog+B2
Fvo1/BEWU9HZLTFfjPB+kJM90D6uepKkHwhljTbBGhUFsFTFtXLQWtExc88JbhRV
Lly/7n61TXSX4ocBhnToWZriAsBjWXF3nqyMYKxzF9O9E3pQ8YM9uMDiV+Ed1B2D
+J938o/01pIVPM7dF7aWgDkGnTdEsoiMoiSA2pVhBSJ+eQwpxftdz5UPFfIPG4uu
pIIprx4777TRWrJ4gi3zwdENGAsPumtXxxw2mSFYItsoT6d2fu10qPG/BRC2RT+g
AzbYOk1Zrls+625KTgwInleyZA6YJiKxTLvoRrvsagpO15bJgxE2QEUntO2+bI+F
mKJtGeYf/QiLrCtGGXBnZiipXvcBQOd2Od/xhH7f9yngVlawfE39wAQduFBjEyEh
sEae4Vp+CJInOcxj1iIYnqJcM0U0Rc+u+uQETv3FzP/f5oG4Ng4SoSI5eNKclVng
1z3A5dpVQKTXEWhhxohVpjywE5KmbfDLw9eyR/sVhJ80WmX9if0Zr826BuqQE3zH
BTPehFxaM+1/9aKt7PCyhcwWuzFPiUHQ/kkQ0LQXiwubBHxJpc7lmzCwuvztCTFI
IRs/hDhTEj4REtE91ea5OhzrUwT9f4nlS1EgYvtGlrNy83fEosNCk4cyh209iCgW
sXj78ueGftH05g6A4fIPU4khac/QTHjwQHv3TxJOjdsyTskBcJ1eU1J0zHreu+4G
ebPhjRC29QR9D+KBKZO6xvYL4YTSlxMejwnRzTqu5DAHElk/5xpiWlseokJI91Dc
/2PCJ6tSyo9kkDGKAyErY6b7V3ZD8gH/D6Ad6u0JWIUOmNvtzqKNA+s5wOjm5OVC
fL5Vil3bt6OKH/WBemuaBW0sp9k/2w+bMOEAV9gnH/h/W81sub0JjM33z1kJptCg
Y2PXMPHR9Pkm6onyQDnFn/5aQ/dEzop5tu2o+xq0HM1SD1H9ajGRpftk0qRScKiv
bS0nopN5neZ5XVSvnH+RV4igLqB+1Rt3mDN4mAWXHg4Q9JGeGIiFis56ZE+kg+8L
U08VvRBMKXPi+Db7SJ1uSh6hKR6A/E0xtB0TuPJF+AsK/y3O37oTS5mgUvGljNzh
YV0mOa4FZtLJJXI+Gn+1jLjMu9hlgsUtGITqVcGaFO9uu2zGQF4gMOOlbdrp0ap5
ZE/1IGxqzVjApdyFSdt/tesJj+dqrxinTgXjhzHEJOFpgJq8+lF9TbOHtodEhdHG
ogevtKtVAw+1PxihhCQ13P87QQGLYQjqzTDbPMOfD0owo7XrlMjLKwQ+geqRL/p8
FvasAYFQpwMqXZ7i3VIPWkAFCb02FcKZFvAhho0UQiikw++xTxwnso5Zs8gMOV+/
iF40dpo80daYZPrWsDckXTbnfSRfgIHica9poO5YD7nEPFggutlDEa5u9ZtAHoUU
rqNPEEgIHwFPbu9kHLft7hlqz9AOiDWK3jhBlLEdtml3hiQRw4d6uqRcXJZt7Ijl
4Zf8XYV4J1KrlBaijKdKmuhHgAejO4nAP4bvtd+YPeT5LdLDjfPnOWiQ9OynNPam
QE/vCXcSyXvVSEVzaEncVAkXKVvaDcy6dmFtu9s6Cexa8tmkw77w03HCL/J/8mTc
r/272Y0UJMoZvUgnD+g157gr7SbjHfWWYXR4CkkpS57/DcHhjHZJco3dEHoCaobm
fcdC/Q22e/jiUZj1/A03EazmBr1xBLlYqS1kHeiMEi1Q49T46FMwxaJwSSHp+LT1
ZHuslYMUAmStue3iOudjYzv0zfaTHqWPo9W++tP37qeAVPJp5BhT5Q/P+P5trNi+
rDNIiSDHKAULprjtp1JhKySbxiTVc1JpYS2ksgI3QUdxfSPHy1mk5fI4fu1u+Lgn
dLoo7dZf6BkQ4puB1aHYp61+HvK1JRcLNcfuGju4EUBtuyIhV7oH+99TbnmwwxnX
R669Ym1vpJLfZigfV47pf50ciADSNw8RJKYDSyz0kOkZG/PP0lExbtxuCCDzqMoX
IvmF/3EkBobbJYx0yj7hUoWhUAPiCGDT6XoxVHaVNKNZzk7p1yT/RZyN3VGPtltl
vAFBmSAtVC0yl/8mytFhln7wTcMUNlQcqDwg1OrKicK35dp2towp62qoy+bdYkHW
NzFHoq3+zMJjJHWBLfnZUanzFXJSDsfc5TeFslCxaGmzeXUftG0E5iClOS5lODtZ
3/DZxXMD/og1b5SA7m8I9UIRhHcDW/NFoZpOWUC1QIWtojf4t1I4uYyI9lV0VAPc
uf9Zfnm0H/GtXl6cUKMpXDe9DeyDRbzwiekjj7K0aYlrDZ6NhB4LR/IBr+Lf9Ypw
6PuFQgdve44f2z89+m8wVNWAbjQKXc+tMcNaMDgjpCgz2TD9Ho9WM4s/PC2vKpw7
sTxwAm5SPik3ern2/BzZU1vOBBr/ZKppr25O6joVqkRgxFnu/yVowuO3XJbXcu1b
Fc0KYYQYV3AO087WVXrXhXQE1KfeUMeJEnVnth6r/OLyUBR6Wk4e1GOxMygOPLM4
gT/CCNJh7Vp/IPFxDt5gYoRQtP0ETqZLdZIhD/MsbVoc7JSgaZKKih2JwJ+T+scD
w5cNix7ANEg4JPzwVP8KAEyuYfo9+RgB0MgL0xk/qaCuA98xQdgdVl3Y4izdB5xs
bT1c2/VtZ6rN9vdzDiDQgL8u9erGrCTCKoJdXkylAv6VDXwj6orXI43pUsG8RQyb
EeK9jLcI0R42EHFwZk+j3cKiwOoavB34loX6H42lpVQZ+8GYEZthSS4oGZtxawjf
/0EMpIfSKsFtMFBGazYYBZ09ChD9mJVkCnDvjQLe/ZgsxFDQrGcIYgJRqQ3vYXbn
KP8GV4XQg/as170BnV9Nkq6Zhaywuz8xZ6CaK/nid9hf57VCZq6pIjjNG0Cl1B0i
rMLqZccmK54Ll/ATX9vsUfllcv9ku2dA+z3/MFL3KulR4aRqck0+1zKaB2KcKqXX
t4/EONdkhXo+dZrynuYyxDdjMcghJnRn6Ujgza7C/gLb62TROTiToa9MLa7ZncZO
tTkVIBfHvvHmBpKDu61wnTROq0/pDMquBXRD9eXntpEU8M2Amv0RbP009lAIjyMR
9NIgiswhyQ41hJnBp1EYEhKe9tvbHI24kz7NuHnxYTtqKiHvY901lt+I9wNbnAlp
tF9bquuhgvQoTYYu5hyKSRSGoSu9WONYr22IvoyAoCuG2X9/DByC6PwqNfFxYNSU
bYqCDEbuJC8Bz9/+eAb/g/w2bq8VWysv9h5cTTWAFmOKyosXbL2lA/PcXDxtexwk
DUVa+VIcqwIzylxrujFsMk0zVb9UiwM8khfHRsenReP2yhYCLRrOyOR6rdnLJEAj
nR6nAyEN9dou3lXPnP3to80h2TzWdjQWMiJtjZieZLIRFeX8R8705Bni/CozTeb+
teg1Dqc1vFWiAHkEG5Mj7uKX3eKBTdFCuznUDDZXmTMpeu7gwC4xgFSzH8oavMSD
0tffLPa808/NAWD68pAMW7LkOsn6i//TSBtTMse3RIQe5NkTrD80t9y2t5W8m+4u
+CF8jpJVuokAz5g/Ex5FuucWubll7+Q0kZEBZoX5Oy290gg3YLV6hQ5Fu7Al7Jkb
53wf+geRRAQ/tHkLV0fQIY6qsNcbhhKMqvQ8uWHGDbxuvWVIATD5enZDFdOpOY/A
b4/7zchTrYYizjSIITnd7XWWFKXPvHs2MBBjOyNeA1q876XgXuKutbn4QGKqmiIj
DuPPvimC8Lr+mw0D0vQ3qtHFrcwkFmaIy6KXtMDEJcljloy/dKnnTzOOGkVyrLJJ
tSOsGwSkHw+c4db2/ejvNEFM+yTrNnSXH58oxKqKeE7UK8ux/6abFAOJpGcFAS6Q
arFgmgnFLpE1F1PvdFwWS8SC3Ys3+SjHBfMSlRKqWSKij03g+LN7uo54P/zr84z3
tuUJ8tEOIGGepa8idq41LclbcntSFrzeH4nEXYp+568TcnNdIsm+FwT7N2vbw6LU
b4ss+9PqHG9QZnc3AwVOku7gB/ZHUM9t9NloTYnJeFMmKicxRURz7X2t+G8TfU4z
03+X1sJzOxQwryiGc7nJPxXMiuKxLpwQMnCTLp5KDJbHzWc/2UVMOlwpsgJylwLA
9yRV8Ka+5l4BR4b8YnmNE8gH8Dy0iLT4RjQvz6AQB51MURbHQN6PQcOdyOzpRVfE
ZMC0O7HhVwIx91gP9l6oI0JVv+9S1mpFhbs8YNk2QRpz0H+pucY5dKjzuhAnw/5+
Q9+U0JBJJN5st6SwUrs5NNIJlpOOTTT5wClDIC7OcqwBz3g50Y+EuNbjlqqQLKZq
Er2+I1vhgu2Vu0cJZr4DUjOAWNoNOgF94vd50WzQL46MtOgGEj+sqx4i/2nUWBac
iWX/alHbWR4neo3r7Euf2GWA2FQUtKC7SWYRBllFjwhW7DpiGrFjIlMOZLuZ3RsD
6b13b7LLYuus5cQXjDxN8CEjEFnKlOnUgCG9BAEgCmEpDDvSvRav5Bs25WYDQz75
co6pBXlE8VnvQb3+wJFiRjcefzdAT6dIy4lZ+z19TCmCZ7X4c2UI58OL9Xo2v/4K
TaTx8MDlOjNqlYTtcd9c/eISSXDZT6SRudaOIIySC9YAI29PXthW/H2LSCq/maOR
HBy/TOYbxbuiIR0HL6h4VtbWmX8UXV+7YxjS7BKPZyKExsfrUXK2LpLm5KQecnmy
c6ZEozcFOpInuKoZx3FQQ/l1Rs4w/mE5MJK1lJ1I1QccUIcLdBB9gXw9T6gDZyud
5S9uzYgI+KAmj/J9Peu7PdOddJigbIxmpeZZy0ZZbHPCMJT3/kxMMXkxs1CUEe5q
nJu6Zt3fBgLiHp6GcIPe7+J9gNmOARVelJZDeuqO99/5rGnvvg9kRcV2ggTmOYqo
MGa1yhUWCH/aQG/yWb5MH9CU4SCNjR2a3qrWFJWupMinOehbiioZpQKpgHbrtRJx
zvQidh5hk7FPwIBmcB0rIkQDKolfc3jjrEcBUbth2m9CQCKxu8xS7PnYthllTRJr
+iOcyO9PoyJW4YfxF5c02N3PUK2n7E/3qlgZl3C1HQjjTNQakalZD9qQeIa/ptD9
NOBGq4w6mashreza59gs2LepgJL0ujY5sAGKV1StXzTTu2bz8fk9xCzJGlW9yPBt
BA48QfD0ZfPLyZYl+dviTX6dhrWZBpT+oK2GkWaDXfdiILQSTV7adsp9eoKWb3DW
DFpnS2Jt0SCifKJddQPLZHrhEvdMbzti2dttN9oJXZDmC3sEkUkZBzmH6l3kQJXx
b7ycgG60de4GqU7MKdZxelFDCL5DUf2ShlAQXeS94TXnoNdHONkGMceE2U82z/f/
74Ct3h+LZc1EVyQtLEdMZ+TfXGlscxSLc1YvBOY2xxhvlS6QPjNBzg2rFOKrJso/
ebhuKEJDqnxd3oVxCbbTgPP30BKvB0tvU+OLk3c5HNsNW4zy38F4T8YrczrepLGc
G0OLR0b4ad/caHA+/91oMXg2qCXaob/2zKbIDNnLI3EEvcySsjH5Vw++Nc8DTY9m
slBg725/Prk53GfkWNDDdLHOKjt6ofTNV7hg5yKqw+rwIPanJpcMjE6JgPTXK6Fk
z9bIB4JVRaI8eABeNJZSO6lzkAQLbM3GZ7f8ZkJ7D5m1SMpAkT+3uJ3JqSog57iw
qrnlTf4veT6yQXeizXLtdxTXBow7cprWn0l5F16XxYWoR9JYSX15KJdIiAP9WKOW
ZBchcM2z6MfMOLrIOONCir2g1Qv6pPsXKyextwN0o6r5+4JOqeeY/ApZ8rYghIzk
G7de8efpIdVPWqnrHpApV7tENRjWvXFxoKciY3a0eykZSLpOW3XqH/oyezdyLKzk
DIJpxHc480hAmGaO/gowRwGPqF4qAHnxQZQURPKieU4KVTdC17sy+hkPiy/Ktgay
zB33Knz9dNr2yQEajsCtgpUa9Z1OZtVSr7t+KXOJp4li/yYzQyDPEQ370dqdojnS
7s/TmFEo/ephaR72w+sPQsOHY2BJ3EX6hIbS2/jeSWeAnOnUfiFxE1fSiS3f8J2o
ucXL2uyd/tsKkZZBuA/LTp/Wp0TbUJuIM6es3b8ZuWwh+fzsvZbn00FeN+8SWEsg
RGxm7p4YJiDU5pr0+8H3gmyae+rrBJP9DMUAq/lTbSpHYDTd2sU25tjWxB+NpjXN
/4n4Epf7/K4Ci3lAXD+1uLbJrNLeQvjQ3XpyCLqOK6EkPEnv0ZCc61A/JJExMZJM
Ihx2vgwxgI1A2Js7s76rYm6MYENczLf2pCN9TxVE4gH/R4WxTSlWF/jt7mKhjNCo
XFPsvy0eGdmoZugRjq39rI7nLbAatg5A/l/ilUEUPddAIgesQFgwUO8dn0HwF58c
7eZvAlkeqUQzB36hPAfsi8txnQIwkrp26PaBnwlpFQddS+ioUH/s+JHMZist76/N
wgFOWORmvf84vmL0sKHJXXAkQdx73J5JYali79UjZhxXk0yM+FhDvelUgGjLgBVw
TsUXnx71UOXhO24ttJvx4Tmy+yhRu63ZtDNPYA5Xs7iK9NBjHg4FeE7W+HLCeGXy
FDZGrty1wTcDHHbIbs1uXXzKZPIVolUyZLdiE6toKNAOF5NQqbPbKpELkD7aqNjE
suX80+nkL376UJl3oH2DdyWAQ79QAqIzMCtuwMX3/+CWK1PVhKxeBCSgB1Asc7tH
42T4mGyk84W6JHaI9Xa1rrBlv1GFL86IudmE90o5T0pmlgL9xvPJZObtab26LfSO
K7oOC6MbBCbabwpRZC8HwKdfbyMIvqRc9gBzHByKPOSD4YFKJZ2+djbaBZMqGLKn
0zSxIsbcr0puPCgeGw6AasMJjyQIs3yx+0dGqYkD1boti8P1TEo1o2GTWl8xWxib
0Yo6FEuQAEinaXSSueG4qYgQTG3xI6ttf+8uIvmscz2P8/bWTC/vCS/Obu1Zd8r2
/F4RMnAdr0JJ3x8XExizDVRebqkLkqSrjvZdjhBPVYPb2BcMQ+Fyi7g8pZVcFoJZ
DqtOvHKeQSsviR7dYcM42qeIRM7K4UcvBzFgUc59imgBIiTVahRyGJTVtOzhuXXa
7F6DlPAXO+DuZbZO8EggOt7EOvuB5soDSWqyYxRQ8928KAEs3usyn8PjBQiEnpsU
32jSEdzDq88hSpsQGeFcnu18Z0DQNgz/2fLiazrHI5LiwIq/J77V32uOEtz9QBF/
VoJrH+fmpo2YwKig8EN23Wwa5TGZjSDwAYbmtFTG4oGifJRjS/Lm/vcsesyg8uGs
8qXMyk0wuoFgW9dRh8pt9Elhjl19svCg99bcIL+BJMQTjsNsTsw/dyu5gz998nmh
/mdjq3VD7yKt9SrIw3pwi10UVjJJQqcft+uxvXMW3yv7Y1xXpgqhBz1fhhPc72rK
1KsdHT8T88GVypW2OQi6/s0XVBg1uSlAHrDj7ylIapKxOwT2qIz9jz0O107Chd+z
wVgN0xHgCNZuEYizgSveY/iUFET9MaGwpyp744NJRMfYWjI5gF8+oRaP3dZMEUtl
Uvzqfg0Tz7WsljyWZ6XXj7xEYmiWC82KR+fN7kz7UYYnv4z3paXhxcDuSd2NtW9E
H9GHV2PUpPP/HrxKdEkYMPAMKeltFKGKQ4urFzA4uwPL36OnAl8TnrADdrOh5Q2X
Q/Sw+R4zsL41bqMiBkmh+Lyxj0rhlu1ga9RKp4buq/a5z1JQBH5wg/j5SxtGgq4W
N1+VE/BMaL9LFqr6tdDN0yk84H1nloPQwjHUPNn+hfuFpEBOexOyC57dQ6uortHv
9mW0bNJ8HGT0Ks5aP7rASAeZuUNztnt0Mwx/fZ0pI4E/2IYfymH+7ErCAz4FXayc
xpLZgXwbX0W/GL3FdsfeG3HZuX7fl8G4NZSkw1xrpDz+IwScZT/ShEgbXNNAu3ja
FzDLTPnxXBNqN1C+f2qIl5yPwEVyskkTQW7Igtb45zOP4B9R7HuWnwZfU/SLYNc3
BwVM2HzE0yiWuRCcnWuHX1tNsi1+jXRdjf66KTWTRkYMfhDfJux/gwxnG40fmz9z
e03E+KzURMHYvFEt/AOfLFDCi5f4EfnA0huZc6REFl5dHNhlDNxlskK6aPHfVg0C
LWn/h7nzSWr5tnc0Lu6ZOcXwdcEGC548kGuH/fueGpTEimIkEEKss/Yh/WowSFli
sylfX0Xr7cIzaLyQnDrsS1fYm3C739PMVdSJ1yXqDgR0eBMxkbOZ+Gndew8wapYa
NVFRaCkSaoo8LYQ1Z8NGrwl43SI0lfF8NPNkKcEGQmnJJoUezVfjbCtyqEV0gePY
tNQGE7/9vSsJG9E5KeEO03BbxCQKubj7nF2XMpmDamcK/6EGxdo7ZpXEa2uNqaDb
A7UNNolF/M6lUzSYJJRd0yQ4NrYG7GjR+R5mLxXPtgfYnpWyR8dVW6tH5YKjRhrf
62GthtWf9EyLa9GXHjiN4hzZK6WvdSNMQXW1fBlyCEzKnox/z2qNNOghKtWbJezI
11NFP1Vh7d/c1QBw1KHzh0UIAqpopjKERGC6bw+ljtsheVmMWdtruks2vyloPnTP
xMew3qEd3biKZ/99qyMdhPQDuGodwhyf/ElSH+C8eRy6gFzxNhLSoue6h+5Uvr/N
UWx0T6QlWlBkxXrhlRR11LSSBkW1MMPN4GD2/Luhs/bUKzNrbES3MyK1gYquZSvB
VN/wd+TFQOwnisxXLDspTgAw3mjbfEgxXldSKCti9fa/jEPqdM0Kc9nEi6NXiTnz
wUxpKb1FmnTixAYqwVKHSDbpZYwWz+r8L7flOg5rj+FeYIYNvbZH8JKMQujLoHIu
QaUScCwlxdU34CZ/jysGEwpOWdSfMPBuw+4OEA5FSJSei1qNZKCSvsh6ZWgfq7P2
W2ErHWNnFzathrAguMB3fAJm0fM4sC2lR9/hspVFuYTEreSWOsHpAjjURfTAHSbA
TeoAzHD80Bi411isIY+LAFDLwYX2AodKYuf7iEOpu/OmPWKOk6PzEtOqhwWE6UG2
qUYDjRgCx2UVLA7w9+yGWmjJs9DjivVNqQCyNnBpU+/wCdIpPtskyZ9hzFT8j1ak
BOFLA1hXy4mAACaqwTnWe62jQ/H50f/JcPeTZWXcAZevZfuNe8EnIKweUArnk1tL
vEDUzovwV5ewfc9OmTLkrO6UcMwNOGneUMoaMhTGLWqUIZd7jFvlICJyeowcZkTZ
4h7c+7DxEA7oIbozTFijBREmK+KRPpyuBF6h+f13nLFN+ahHfUn4CtFh7C0ie5Lt
SNQq/LZXvvIWz+zQro4P7EcmjB8x/WR4QCqsQnDqY14X3lRv+owDk1fbbvnlCRXU
uQ+kH07R65/OR8/7YZfl3DlA7tLkoBdtwoi1h9n6/UtvXt2NrvalApjlASEKzoQS
ckREgJgaNJfyH79jhoAiSf8tSfUJhw/EWhNdXVKDn1ObuefblWqOvwFLnqnQkA+S
NCdVJG0LXAdOlJL4v1fBU17njbYuaHStol9YheIUttZGkw4qnb+6aZCZV7ORdkYo
/hx4Daf6TyA72FEWunBia0R8j+TTwtYFA4d1oAHmW6HYt/f22uMWwh0Mf/YrxeUk
1gcXA62UBLvqzrgkxTgNGqsBBEFJZZz4laqYy9fxh02VTHq7B80T9ZjIvwR29A8+
nNB62rsgtQT1zL0bN/fAbsuN/y45vhKyBgcsrGVCvFZo68YwF91OEwBdz43CxzDx
xICr0E51nMGVyGPCgI0Wj+ewy3+sBlA6D26Cydq+fZijMQ0rGIVuggPKD4/XuHQU
i+Z7sR5eibleCPDBD0qW3L94B2oPc90PtjCLZq2rpxVmPqNx71Mlk39/U2ha4QKP
szSqedgUMiKwmD8rSR/hSXmVVdQoSaCpI8Fu3Sqx0ZqFuMne+Gnk+LQhoS03aPaq
j9oAwr6HiqD9ZmMrISeMFjUj0JO7UuU+Da4mUpk827jNUvNv+Jqz69eFyTAJCJ/W
Bw4pzxsdM636rj8fOg96QTD6xItIRtnMKIBxXX8IQx+HNE+tpYW8+t8Bn7zlwlEQ
Lyps1M1tDbSvHHjk0xv81aIfWokhkCUld/eKf05STsG+J6XA9n0uJ2MS+jnc6Dnz
JyA4lFJkD3Fj6t5ao1HSwi4l5hsjsWWARxRjWyXMi1nHWUY6qmJ2+wBaeDoqZR8g
IxVtDkxUYMWxh01DDJyjvws+fZ8BZ09moENJ3dLn38H2a71mXdhveYhL78tMGUNI
jEgNc33d1Lc8tVIM/EJyBAwD4yDrAQvkYRxSs+tpGMDuE4U2hRl0qvxWtCn2OOJS
sE5j311NqvX8eg6NbdufhS+/eUBYPyBax/xzpeDQB5hdHSxQueaX+lE8fjiFtwkQ
unhjEQnJ5J9utM4oP5XQLNAUeWRa7j6i1p9eLCpFmLspaYwImEl6bIEC82Rd+bro
1LO5m1LP4dufcl7G3wjUEU5sT4HPvEWYYAdDJ28Bd2uvJVRiwFySHcUe6pI1SOc/
IIvCRKFi8i1aWzXjTAg7p84uPzK7fOyrzhdInDl8G0zqwpPmqZuccJSzQBoEEvV6
cpqxCK/XQmJ/Z/V2hiMfRaAjELqEu9JgQ8SvV0fv78hJo87N8RN8DIMsTNCPpqaW
cR+jtb2OwtuPImWfK2X5DeMatpUPGMDIGNSpyUfOyzgzRWEi/SBhWMjYs0Lf/HLt
7hlTUqsaMDlh4Cyzt04rx8krGrMw2ZmJLFS+it1tO3xbVvMIAP4qwCa2YRUtclHs
Mu7dq2LyJrdHK1P6AK7vayZFsKZpzJc1ylzrmxZLppgnlSOaAHNWefctzPUw8Wan
xmakuVElTBAfMQ+xwSrrSmfl2xQeoqbWV5ceDj4K1IGw9S8YDoY1dGGcaX/PXj6M
pc1Fwfa8m0rd/nXXloz+mYXNV9U+mV9B9dQnnhXiIpSVzgP/5B4p9qRrhY7VxrCJ
EcQz4x23iMnX5Oj/X+dxYQFq44VxWp/SvU4X+tlpYCocGrX7Ml0cUBmGeS4YaW71
DreRyAFVv1LYEfvA2AxgnnlbeZEwFZ03PKfs27xAU6Ap7UsbopWJ5kyOIH7C4wa0
BggwY1PvxQVVVat514pDzjru+Ymm4OYrdlTBmqohLPGzqXabeUeu1ydE5XDiDKZJ
WmbM2H6D/BJfb7XMqXWd62ooGQnsJTEF9OvGpy1+YdlKSn9BK/3Hp1GIffWQuhWd
JyaNPYcPifeqF/lchu2WKmv1N4SuBRrhtWw3sbGJvlpecCfQ49uYnUZLT5PTCgVj
ZLdXKoKxRuV6B7crlX0hb0cBHURdN7VzKHjGPyP+x/hQyO3yESzWqrDX/I4fBZx9
bGkYjgSwRADdKFAKf+HhgPuNtKffynxEVw3WmCfBGjrXgm/U31gDepzyaedEydIb
cJQqCCu6CPTVQ/h+ZEJu6eNs+1KcUS3q11XSYyLo8ox/AWKLdYgIb5F9lqtWrK+e
pnoeyt22Dy/maqJxlGbdkMZtUWMa5oh20g0SzJoPqe6l//LIxkamXdVS7x7+3kYa
BXo0MnV0SE9i83KwfjLODrASxEhfRLByLbQucoid3rCJDWdubCXJ/TkYeQb4ZSiM
+8trS59vytIjf8hN74osiAA2fqmtb3XWZ6561xyWyxcaLdTGzZqgVL+dqqXy2h1u
S2ucSBv7dspAM+RhHwO1ObI8tLwvlsvmY8uZ69sIFhy+SmpKQbIlJe+fWMo87ZDE
iLmsJ+8n4tg5kjqa3DtBlN4QDUsKBDDpPTya61POYLsMBZvZ9iE9C+FUef9sBv6v
YWLv6LqC8xgh3LUGWLQpSgvvUBrd6wt0Hoh4ocexjYUG+FgmdB5Ca+16ZH//owjx
fNOl1sUV0xOrMjk7Dp1PNj8uxCBP27aOj1rxeAqeI52hJKsMAOmyK/UZTNh7ClIL
8rMGdZepXDrTPcxvVIChutfs3yp3FUEVUZVXPcMF7+hI6+FmDJeY70st8IFdMtlC
NlQJ3wTAZvRIvgS2LY80nCF5gJFcZb2JaFmt9t30NMgvhNymT59xjlqK3nT4NO4a
6xsniTlukZm4s7OTtMfespnA4KfSy2vuLr+UWGncwrFQ0ME72PSNs5vBiM8wYRNA
6zfT1DGKgtSGpdCW9TkRp1/XnjgHwhDqeTsbxeJQpv0cxsS19jN1ysw+fkFXaXWv
CklZM4XafyEg8jCFX9FDf/LpQJsKBRFbhcfXHcHQFymN2jXgVK6sPVLXPL4p3mYg
+HSJcF0LBIZPjG2p9QlRlMtGilXLGev7ySglzpCbcxmJzShrxlG4ZpYKgnw1Fb++
yt8gi0ConZWB1gXQMmpe4Q6BSCXTwaXaCRU8D3lPgzLjCPj7hYWTXFFI4S4HkfIn
jgTyLGBHGnDIoEeAsG8DCF6e+PY5Gj+hxG8wzAbxBgIa642ftl2LCorhoVhtmG2u
gy1Olt3bAbjv9u5s7berFOu52cVKt9P5wkPF7AmpQoAKQZX7CAIPGKwhYI8sgV8w
uFtBo4AWUpPGbvO7UdBTfYQKs1W2ctSpLBXuthvwt2VXgp+DRrF0ajR8DbtjmOJE
QO6LsUKb2aXc/oChGmylpKIHvFoPCrHJZFwDzjMgeTvH/CAgPCUXG9V0NTGyXsWX
gju4TrzH3883O9RGF48vhE8n3VQ80mi3Vv6IxzRbLjtgJA+mjfNHX8fu+dBBtJ35
+8uug5HnE2acYPo9pjIH67RkrTXrj0Mdv68Y/1bLA2mbicppnvPCVIpVWCZJDdr+
Vcp+tch4BcDlRp9kXlqxdSckP5+AuonBEGlsZnFssO49uCzqZQ51Eb9h/skrygrw
LD3LAsdqvrazd9HOLW9UdjxP/Kj1N2bYkuXEch0JPIRGk4D11q+tpCiE+Yc3LI6s
kkc22/d2Z8s5kfj3VDf3ypLW3GpaiS06XqsA0YM2MB/zTpjBBgwaJUueHEMkIQfQ
m9BE9ZYQ31uzOCCFjYVy+3C12PvJgdlfrKdBvguTTw7q9Feoq72naln6gST0i7zP
Eo82owzi+xdQGwnJwh8jKvvisYNc2kfZJH71fQqbAc0Lq1WHv9r6kYk//8ewHMFV
4KdWWCeWBKR9TyYfLRxYviSF+hT10L0+I8Dbug0fEF4+E4r2mcpR0WAk5YBNBUm4
esm8HWfzubqqAo61ZpGI75K8za0fsjoZwzxESbbyzaRVsSi/nFIM0AZatev2oy8Z
Ju08NILWAAHE4WuXigAplGAcTSA/qMJyn4Q79HLXZLg9qAVik3GwfWpbYYZRaMir
4Z1WtoLNK7nvoi4lEJhHtO+d/x7KOZr9l1RUBzLqho9UZPz7C0kFStre0N+01ntV
HC9cSpWy/JoyCLJw72RvPgnSiMKdzsOgnKqPKZvFea2Adqh4CslBeaDYjXy2+5Bn
tPfCU7cvYtob7M0hDI79pOIQo2ROYZfsyQo4U/28Vjgh2apgWT5pBQxqsM5f27xD
jgV9k9E3fgQ+iTXIoreHVthwtVrmN1BSLS/7ZcN2fW7XEG3RZX0N0DRt8syog5q1
3+enJNQkrYMWk2nT/tw1efJ2C+ckpN3Jl9Mcgv2sxthWyr+EWNplfanHoFftmMlL
6eR7WrvrP0PhUoXaQg60RAi+4BizfKxCbihIYukYaCX+2mCEstVWGm8W+x016EUk
IIgTh3O1xUC/kso99cQlolzQXtjfaQIeri4BRwG7zCMkGLMPy5iqXVTogFU4Ikuz
MSA3FcciveWsB+SdcYPSBWntowPaORsnlmFBWhyHeJpByl1a8vx2j4Fd3h6aSott
1b0PMRlkcx6AitVs5oSSU3d0pSB8dtDEdvPlJ2Itcbl+M18qSUS7r1kUNtC+VgAP
u9R4eOBZ8Yvrb/4ks+LObKVPqP8Ua0jiTy7jcQmMoz4+SAoYiUe9RWY0AHd2BZuZ
rxoKI7yIB3W/dajpq+txjzIoBj5uZMTKaZOgOpR7q049WTBaABz7HXSm7Y9SCZGp
AgbwPOz1o+5P2eIO7lHAnN1a4rccbSqQKruw32AKf20XR0mQx3zV+hh1gfVLaeq0
/L92u4cpqi4NfDuKupcs9kx86rBQqclqExhzmQXBUwtKQY72Fn1sYZQhGcSoDmQV
Xy11sgcURe3+Oi2FzctCI/Be0W/eTnCYocvllXO66M15JzsnrtN1UuShx1Grg1EF
LmVaW4SHJdSaZcTvqMQggl1a2X3Z8x/jakVMrymn0868hjgTSslksnfianiDjK7C
RcV7kYDnrkiZ2BmGoy+w5OwiJG/mdW2niuSYkl5Ewbt9UBCnHkl9a74ScyiZovN4
H48l/ZtSp9Qfwphm1bFw0a009BJGYCOvCeT3DJ4usDlfkASGyN/rwfuRtVznibA9
ggU4ZsDKDVflVEvbcCa/+ohdOc0M6goC5cYsyDOVJ7jNGmmZxQDwDQHoRYknIGCn
3jocWtsXrTGyMXc8a/D7dXh4hmojOrlwLwFKFFc7Nqf7bIyE0G5ZtnFCTYFny+uC
ivmRMUZOs9FUkVfKYqAJ2r/WJ0WUaWnJsDHybqR07ogzIHv9ZhulCU1dw3AV85Gq
2XaB5Z8Mx+bQ7u/ODLM0xCA2GyWfAbPs/EHzMDfxyV8BZwcZPQaKR2z6PWg4UGvc
2JA3FKq+lpOyaxEEraqUbymlU0zvmVUKGdlDtFprpL28jMRYZ5K84fkjMlLUZINH
hY58tgSX6IWpF1nQrzL5P/HAPqPOVYF1bm0LqmNy6B28C9TJlEMo/7xm6poQ0hcV
b71DjWIyLL+yNWs2pWSq4i1vQ3XSsg/CSASTkP5JLDAPICzy78p/sxpYIxONv8/+
1GAtGp/Bh0UhVl4CtQMxR/rhbhpkOOs+gEy4ivLJ708N8zOeNDCVT4nsPaP4GzFL
GBv2kmv/Lzy2jWTCc1N+Vx/oSjRIGUUfs/7KtGux76ZaulRIYXLKV4MLM+Gcx15H
v9UBDyca58E5X6aZDCW+OiXXMnemBzvGfF7u/StBZkV4etSdx6zwM6ANuRrAy2I9
aQTVrwubM5NSXW2/RLBadb5DD4pytMmDy/UAS6RxcAQ75WxLdYjeYcQljZHoDCTM
MngMBirwP6WC2YI+epBXyiq+pbqegysrk2+Y6zxSQB4aHwc98YmHGXVbcSftTDza
+u2pSKl8OaW/PfhksRgnpjfl8zofZBEniI3Br45H0huo9o4yLwAsXc7PgefQZvWC
jG2g37ID3FEO6OTdDG7aFm+fZu7TLunFqWOiUVofV9Xe3REG0bUjYisENHXP85Yc
9kP1LyFnH3PciPOLE3VcTDbTBzi4OQChHyoFZ4lp1DU1kwE8MaTrzBgpLgU5YrfZ
XpwBtb+YyxdO/RJjQvY+dy8gzk67swC/vBwi0uwSIvkJSLegGYq9bJELjqU4+B+n
/VxWIVX6Mra7+31yIihMvt8Hat4AK2/K0EkEX7ccjuZlk5lCdisNgGTFisO7fRTX
FBvDVehMVy7xu0iMqHR0qAd6iYwu1DbZrLpx+fL1RvkB8vtxS09+iTVI0LnhX+6W
r9hYJYgjF4+Tb1Z3u4HbdgdR8GdQozG+Gv8Wk5xLpMLSV20sX9acajOoVruep/kW
b/Hv887U3hUPL3BkmjT2V9KpdMDk8WjCXERYav+Tj6SyZhX0IuADkF8FJHGGBNCn
YNEekPq0j7UzXwZtfUOWATK+4ao0G0w3Qa3QudHdc6wYihqeujmldtCmmp8Rjkz1
rfMtzp9a5n5PCjQuGoG9l6XnOt8SsW8nsDM8V7yBz4GWNrZtRymaPlrXd36Fdjd/
1FjFGydxgJfsuiiEVxexvUY2ZAtlB0bMfOBqlhPHoGWiJzFJhnYpemjIFmzyYUos
+837Ib3nCoXG07Ebp9KgegGsc/BJEHsNfxpmRThSEAcVkSRLGTMiBcm/d0t4pUmA
JSwe5L/IhsKEEucyCZs46sPcFMWKPJ3F6W3sWrUClNMtakhzWNZzHpzZSOijCB+4
Z8X8BRoln111JFDH2FtQH1U0d98AIzKzrd7YprnlweVTAja2q/7Nu95YPVIw4pEd
Xl4DAWGMu4V9w+xqxiyfSDY7SRsVkbwcQ9CVDuDx6Uk9oS03e1YV6wgy7uS0wWvN
p3TY+BWNYpTW53yG7b0N5TNaKu0YNOgqR0tL4GWjHTmwat+43e7UzvWA9jDaq0X2
eEjFKwKw70TRLjSb2nwV1tsPg7QUtlIANsZTyTffNII7ajWktpJMByjtwTIBy8AF
WHXBIHKHeS7x4a+VugyAlx4WDkXG3WQvDBp4beLxLmAKoVTFNkWLl6PsnTcukqXd
gavLYIxVD58UeE1nRylWjfS8RyTIP5cMo+O5s3f25xdMZbawHebb9A078Qrw+xhB
oMRsuv94ppZ8NT98CnUA96J0iC7Ycl7rX2ZWyo+KU6/OA+vmiEB1OtnZtpii3Vou
jzBfuVI/k+V6pCYbhwVNlfFRuFrlVXtyO7sMfZRpp8lc5QUgOts7g+mZp+NW/r0a
aMOvvzaA6/ek4wUjxV6J7yIt7vTWjpezcX0p/7YGnZh7vFMrgdy4Oi+Tf5FY6abn
kBXZMSQa/cNfLs/fzAfLX8bR/iPQwui2MZB+O/11LOJPm5oY8vuql95dROMDo0eg
M8s9AimkSVJc7VRHAgdlYvRlLU1IiSkyhHuuhuZ/XwXIicg19q6e1FMjBfznVlvG
PxKIbCMEc8n6WGqAU0aNgaFjdXyZ4UEdoeWfjx+rCQ5M5xQK2VAHzMDUwUlJPNcc
9Sld3uEPaaQ/WATXO1cqpPdJJOuY0EGYs/7zXdqXNrFQ4Q800tBRQZMDIoA1lZeE
Jdm8iaeSCKZpC2kTRhUu4sd7e76Jt+KSvvh2b0pJwYgJVKLMVlbXfYusa9pGwIql
ufzCaiaicw7zdh7R4I9Yus1cUZSiC2HUJlQWH+RF/Um+yIDDaHmjJE6cUPGOBDAs
hRbdC816xfoq9+lzYNv21XS2Q4SRgoQNaMumyCSX1yv+Nda8kZjNcyQdnAL3Ubd/
qYLcPIou2W8N/Q8EIChfwwjD0Ga84YAjHXeyu8jAabWczc5U1Lqo0VjYwcQkePb6
6zgjoO8Aqv1puOveVEOVZ4AllyIYrUh2Uik4Ags87VEYQl6QlGcPI7aahx/+b8p7
R0lXwX56YX5jLNdfGVVQ2XV3GT9+wX9LTe2Zx31fzAe36GMVkdp2a++AwQ78EEP4
DKqJ2EvYq7g+JrJXOnvGzDGCBSzHnPTFwEuwYoELNtKuKFZvo+K/R8+UzU5/EDPJ
I8/ynfI8JL938RTv2Gu6/bLcGuaEm0NMMu+e2PsOrgE0AGpTxz7iOxp+zR8hUX9d
DODn0pj2rkfjCSIri79ID3s/GVPf1OtiTfAf+5BFwiO6edV/b19PUGNk8tuEpoIp
kiw1WhTqNzbrvDrvTzLKDgZ0U9gP2DJwjk/SBk6ft4YbZYfKc4qDF0zVl6rk7kqJ
FQcBohb3wf14g28wP/O+I/Le86Vna1qlyGX7qnHOq5+h76FpoMYfxYL7lr7k4sJU
l5dy+Lx/3t7Pu9HauIi+wLj6PyMgmRh1JgyglKiYhnFmWHeRVxfcWdUKlsL26HcV
9npr6EZY8lIT6XVAEcjxjf5tcXoO7ExXID1o7eDxI8/SoRIZfQKpM8BrNi9vsx6N
elc/TzTGFIJ22QVWpjRAoSfskoUF6vngHlrTQ41mCnZaFE/3jw3j1bB74cyNfwLc
uQMl9X6cEdb5nDRdyHku/WtXUhLcCUpUNUAlPOU6/KJxaLGYdihvKFrDsiSvprsC
TraPHXp5Dv9ONEL+7sl1coOcQVAVW1PluZWaFIG1E0hSsL2SsaHM4d2kpy/tqotp
2lJPZN0aGCPE6T4Sd3Af1/OTELkp5cm6kvfVUL+3Qrjv4pp8l9EnJFCJNdy1YZGs
j/5EoXEkKP1Hvopw08EKMbp2gJ8ah++OL+AqCfSH1McGZVHDjViAZUKcc+ID89XV
e0lHo0xBxrovVGIMXUqPrl0jxOwjrLI9VfnHWNHtNbh+swVSyP6g7dWAIKDIAJkE
PT7HrR40Os6wt23VBKBXnyuVczHL9EJgmaKUAu7xHn21XmVB6TOOWk8BnEUMwQsj
BwF0UOoPZSY7/J7lFyS12d6K788ZLo6OYlBKXJofwq0wqAet0+aBJbfV+NytDRqe
qdLCDo73VHDtCFkOLWWMn3qzlfeiqvaw1kJup2e1LPdNom45P3xDi0u5GhS3lppE
VROLsuR9NDIit+9hskZooXK0g8NXbliNO+OPcdUrT2IgRcvV5o9B9VtRoH/TJkAB
nkGDZmrxf9vqVWU3oZY9GgfrmCm25QECfPzMpIU2cSZaU8B+9EoGFGzf/z150nx7
RqncQh0VB0dP6kdAhCT+Hp2aTCRdkQcTDZ+hw0ibM8ZSGRBa1HaA1XuW1jg5qiyG
g7kj30oesYNtk9Jd4iQ+AT92fA7NdMHFQbsTeK/xzjuyEto+N46vnipO1bWOD9qk
+QcpGi/Nudvp03jSMDd0EXK5Z13mvwwPd7lR5GvoKFfzJ2Qyqu8AtKb42Tyeo3Hl
iwTpEDA2beI+FlQel+dMbZla9zRuCxPxLf5VSIdxQ8NzDMLRk8vv8/P3MjqpL4r1
1bGYROyKhzKnfOley1M2odoBO48ut8YFiF08YTcQvc8uoSr+S4WoEPLvfwGVjS2/
eqqcto3zCkEF2zXHsBaigCnKiBvfi2XJjpfsWYigzKYCvqAYhAhNiDyh0StbbHvQ
oHOfraAUU5+RbnvPD7dQzqXzRC9WGAPqVPK4G50IBTlJDhLPhwNA3RIa3OR4pDWR
dpxFpMVR+7VVEd9ZnX/nGdJFpNiHmFgIXyvMxYOUxAL5K3y7BRRo62FmrW8oHuIR
87Vh5Si6LD38mU53D15nURtyi3ZdS8tJcinJ9o4qKKjhwkcbrQHpKR2s4KuihAHL
OqrWR5z9ORzk5FXMCUYmD1UbmhRDHzuLWWRczHQY8eNriFHD+rp3Ez7TL+d7tbOo
pHqXMLNhWHNZLZaUNn10l6fEie/IWu6ciUFiXe1FahGGZRoDqOL3dT9ZSWyqtkEW
Lbu4kLBsXX/4WNnFPIIh96iYi/OmWwR+xSXe/R/UTjI7BleZzBYA3GRmHoH6Vm2p
vzdWUi2VUxU34CRU0P4tbPfy4oSZ8Ix7BBY0letMnSs6Xgx+HRG2/umdqTXVa9pO
UKA0m0mbdahwT8luQMQBcfExJ+nlRdDDbCepDVOeAlnJjH1YozFl2RKelOdIlH5T
z7zmV8Qtdt6OK6IqXectzMp/vWX5Sb96/G6SKwQNlKJO1JF5TNyJ2+fZyZQJ724n
Cx9MusClYGwFZVvCgHo0OUVCftdcZgap7ATCnxHiGEf3Jz+OL79IDzx8fv+heu9U
qL2/DlWxpyWQdfbPkIrlAI7s0JXbaRxMqDJDiVeSZD20F22WHXLgBVvkRCW3PEVn
70FPMYn55Cpf82juYD4uTBaGc9sE47iyelqVasLWkYX7UIlskYLUSCSA8SD1GbgF
vwcgW5Ql5Yd8vA7SsQoXsrzJPFHidIimAHu2XFA+LfVBxqMVh+27x0lrKgtgpONe
Iz8F27nHATiALV3Qf1vdyZ94SGJcKQGrGZvH+c2WZX2ZsCoSxLhxLZ3htqEa95TM
QlbzcNqcclioW620RIGduEbTZBZ4gNxri38uxzhk3OOiPsnhF9K99cntiPKTSld9
bbFyIbbhBl9h40zN6c0chKnkZ6A7oaNEaJ3vuzXpIx+urKkB4iDiMP7RltQg8qCG
v623On4Mohe/lzunnvKFueypUgCFenJbtKLt0ntvnspdQRC2ddJz86SbC6ML2IAh
bjt0OOIevptBQRsoN3kU0ebFoC8OHZnSCLYgnE05eAKPOcr0TZryMU11W2lbe7on
WcdPaJCDNwcbXZmdf1YJAmREA/NIncEYSdY/bry8ItjUP93hBb76LgL17FmHv306
fOvTmAQigUmWRKmzFnXGG9Vf3nw0EQwd7zcdDlQd5KILCO16IR/fu8Uk6eO/2Npx
szAx05gVyWgGw3ebF2H4FiOVydDHWgosNGgAkq9Jclyp3s7FkwF70+597F+yC5zn
wJxo1bD8KV2e+s88+Z37A2xA3wuECYGXhldrqjFBsIu2DjhdpaeNUpPNPmrI7853
gI0WHdqbu3xBzrhLaYCFc9cLpsF1U6h8NWC3cMBq0IvfKAFg0n9EPdGcxXTbp2dk
BI1vM02/1sIs0ey+692fhgU/ZJY+ZitKDz7wezErGbL/Lad1+bcf52s5VOJi8/Fi
Tk2m8blSX+cunalxP9D1Uya+q9r4tSQ9WHYk+81ZoeP3Oa5iEwiOCodRhbIXP7Z0
ap0jPE1+wmUePGenK3cAY4e+cPu9+hzgAy3FzFKGgWsKHjczIad8fBIHRojOe3ES
PlkmhiCNcQGtldxRRa3TmuQXLoR82lxSRLg3OMLt5CCdmX4VpXjjFrEUBrotvkCO
DczRItx2QkCRftRgnBQ4AhfQnilR7kZS4x01mDpdElVBrUSI48l0CtOgnv290Vbm
iqbpjUDiyfJO8uh/OvXQZTzalDxVkrSNnn6jEYLqqbmWzOEiLbPZD3NiK6o6ddPe
WHdCpjk5oy2lPGJkZHOEyvF6+Gphg2VrpYNdMNbnoigFdsKpt0FyxLp5vNbG5TZ1
FO+gQoImSHJE27qw1FQfT11VCgdi6N43y+0FAkla5MmAv9R+pgePvCk4Ck4LJt1J
jQPaL3gTs05ywcpgsfujPKekpGQ4KB6DzuwgVkPjDfnFP/XHJsTfbnmZnU26LJg2
q7kjeHR0ZFlhrCqFxRSQg2pY0hvosZVeY7GLWFy8IH+ZHnqYlzl9/3G7qFEG4MU/
ey2Ra7zEwJh/3ISV3risSnxkRWjiP+q8Yn8qMF6txopQFxGnHSBpiOUFDFMk3UK1
HxRg3rnDKPNlRi0jVv9PVuPceuTQc7+G1uBjl+bsICTq6b31iSL9u5dzrP16yjan
B39qMZpr4NKTtzA/AOjy7cCXl2nVuj5RhM8cJxbSgsyGB52RaZRZNShx03GKsPl0
H+PHjomHaa1XPwtnErhyix/sM5zRxA3IaL9hWK9Ng/M5+4lcvev28/LxRaqFlHaM
wRUj5wiDy00NhGE9deehQm6h0n/qKqRocI7wPjZbhhlduYLN6hhV95QxkkSCviyw
+RiRYDmIvkBDcPk3OUXsWa5gueK6J8EO7KtSpJ+RJFGAnLeqhVHw3uAmCQTfRkGj
q3puYIwzXFHddgKAxu3Q/xQGAUjZ0Vn4peSKphUfN071HOUr6XK+OKh74kuZnC28
xQCu/5OschE5cSnC6c/p9yucimVUCfoLnoteo2sjuQtP8TahXTGW2kD1xSmpdZDA
H3B0Wp7taKssiaG+WaPsv265FJ1FaCgKjFmJK1U7FTeVmow4jb89UrKJWL9dPIHY
0ZpwYPD8693w9MndeXopgzVfbjPyzQxC40Fq81WKfz5m5/ipBZKu3ZnxMgXqNPCf
OBV8QHNmdgvCCUKm1KNpi2eNJEmxcC5LlXOFa2RFThPjRDbAFbSZp5W1qpzIjqEc
i/OJCZh3NN2ghhRZyHyO6jIuCYCbVj3Rt6Qlg/xn57e2VW8y7qUFZl7vxwxnylwn
1ztJtYBJKDZISP4kb2cNJoNr091I4gqClRfw1gIMXMcBYwSSYfF/LUHF+N0HDjG0
Th6m5vJlCOI9tvmpfWZpQLZV/AKN8ihf/7WzZeo2++WKZdYMU3Mcw8HEMa8GFB1I
65JtFRd+62npAr0wfMPmZ6gXhT6rec/PlREbffYfBGL50Jk/n6RX0GRnje8ZH31q
elzHaE/IYkiFtJN61wR37rey8Ey/y7f8zAD5EiKGObhT/MBYhBK/Oga1MvUDyw5Q
C5enCKY5EV7KJ7xa46f1OzaXRyhnph1dXWj88Fb6pXqaLNbc5mF0djZqWhn4tkAB
ms/JdlN8L+DU4uzrIvNyb1ZoFuByaHHPv28b6OuFgoDEI577BIibMmII39qg1X48
hOjKiXn8QmOuUSq8onZ0tZbh/glxqmjAh7omoFwzuqsZ63wTC1JNWGVxXsoTSsxu
tCQhLaQRaJhZ53D9f56UoK1ucKnZs9b8zAdylmbIg4hlUXnSUjgtGhjzEoQJ0DXs
CNKiGE0PFICLMDfNBtkc++7tD0YfvTkoLsOjo4yoq0oFNUaZBRT00XEoUpiJ8SYu
BYyN3rRdszJXZmLXJj1qEqUvlGh+UK3qaDlaC+X8Hv4zAc2XTdHrGpxl8Zqo/B9C
FK6OWcHjf/JxFKmMHOmb7IDns9yswm1M/WBW/KnJ4d7XhTPPxCBCl5YHJX29aWSW
PmAEW/+MLJLl56C4ySjKnav6jPYcCwlzer+F9kH7h16YXINdZ26BAGGuC/+PjnG7
vTRCbjN5uXV6EzkVTWoKas6oFM90vZf3W027Q/RCXzOv+/DrOEpfzEUy33ny5hAE
abt0TpGSMeW3upmI1OBah+WaTIWEQq2czXjW46guA3HUXnnUmaVqFVIZ5vL11GZ/
BD5Z3glDtI97ulmB8kmzThee6gL9t1qKY0X/vSdCgOn5y/3hP2h6Wym6xot0qrGR
5p+Jw6erzt4frQrqjXImEtmgEoj0BkGXpE+aNRLnpVCjvtYMFu1Dm98upo8Wm/oy
ZzaL6YMKfxsXx/kMzT3K56Kvvt2mFwLP4qiWtDX/278YP0O3JLEq7rT9wWGIByOE
AJCPYd6sdwEDrW6A9vF9dM1a6le3ERDdTnFaiVEHgnqndVh8ynQcENQ9Yx2H6iJ7
XuQo/ft57vHOEPnL+8lE2/d8D3ReZPxUxnFJTeGJodtBUUR7vXE1gQHUbWQaxxAb
89anEthPCIvdK747XUg/XhZtd09HODniD/aki6A7yLTA8Yo8oU8buEA00gq8iADm
evJkdQaqQfQogHaHQFtKkOhR+aKjiW6fDxVgUCSwuJlc4IRwTmyjA/Sv7UkpPFAV
e4Qcb2D6NZc3bGHAKcuonQYLXSK7uMrQ79RcQpf+SS7VdeRNJYgJSpKQcipQVRUD
m+Ew7EhpX9eRvIA5Wy85Gp7JLfyrwzk9dgSeeqOiGO7yF784XZvtorhXMliDk0T1
7gDrb2FFt9fqpixKyjE0jNTbcf20zfMk17CoK4RsOf8xD5YMXMPA4MNL3VuBQ53b
cJ7gTHhzo2GlPIbT47nTKeKCA0XZz/xvmpvlJHSZlc1bsR07yt0aTan/kMqSvN6R
ThJpacO6Ng+P97KiggAmQbwfJGP5oI4Ala8+4wGJoA+8buvRvTxYtIJGghBjg6wz
Q4SkN1EoWy9XewiYwCQz6QgKaPw9e/+OORke4kHMDcKAE3nero8DDoi569XzqYs/
aqKAVZ8MF+XRcAQBQ8aT79+5/FtDLuZSOec7Ipl8/5o8EtM+/UdH99d/9plRO7XY
iXqchVRnZzgduEf0S1PKb45wd34p9ihMZwgbPaz4Bt0a20ZfEOcCYMy0eAiaRdiX
hhl7GLs4rFVMA93srbRtRmMYmpJwFv/4bCWEd6K17iMsNHLUSC17a0NGmvWD9VRG
a5PHE/h2uHCR2jghuVhTOqH04+WyAdba3qkEpVTnO0gXYGOvyZQ+eCYeqewobHGG
73cjyAwn/UMKbdWrxPQwz4DbNbmeHOQOGniRImCU6x8YUE7fRHDaCkVo0hB2VU2A
nnoujIi08K81EJKOdLk1runIBcwtSzviXFsqYaaKFlfrdm3i0vp65od3arau6Hrh
LcJC/FnZ2Fht8YoFDIa+AkgM3EobCHdRuxq+ClG8GTPXpwPdLf9oTFvbxYivGwgo
k1Ei4gnekjtDmJjWdoFBFXbBsChDYoVHYUJrSDTLyeL2HEsZZ3D8inGCyrNU/5x1
JQ27bQADT2AETn3QR0dNYz4sKn5FAgWlXAMTBBfk5t1NGB54CK+zER+63SeiCozB
+1RsXP3ciBea/hEvN8R/6IpXhraJ4ZEtdF0b4jYO4Eb18eA9EirevdXWKwVKIntI
FqiH5gAGP00V6Ae1TpPkje6dAHGpWq3jy3cwQZ0TgNs3YpyBisli9vjSBuzQxSfS
4sWBTU7STUB05kZwuY51iMloNPLH20p+RtlQw0U9HkOJzvc/W7gaezAbFbRGAX4O
0PdghU26tVZOw2+Qt2yxRzC2uduxmI26bSRM/RfyKk3+26heoCC2z+tNmoFr2RDz
wanwE2947NK8xQ4QRvu6AMCuCRe+ZW6XRfRIA9KXZBp7Fq4oYRmEm/1BGg98gUpT
PI88Jhuow6soITAxQLp26I2Tx/KRM2uPhOkSYWKuJhsrB+vZQTpeZp5BL+ywZENI
OYlZi/wsE9HvTsMqxhhUFyjzZz9QkMMwLeEO/ZIYIWgDx8GQD32FLzLjh69wbN6Y
by1Wu6yfk8Q7qUrZMFXwD6cbOEfJtK1MLfRD6YusNh0HO2tnDp9l8q98wapCEOJh
dpYQDOKeyzCU3/Z4Mp8NOiA+Qfxnlsf2uYiyoWoEBeMgiOad0c9d9VzQMjlpGSVF
h2eXwuEERitFvz64n8OwAnTGz1LpJjWAJwmrAxoGyaAvoaAZOFcTY/Hr9309Zajp
tHXvTYSkQz/UiWk1QxpBfUf/jl3gF0Er1greJ2FElwLgI2oWIq/A+m0ygA7zAdar
Qn17srmR3sMm95Y6Mbl00ZyoLZQ6owCZ9wT7fydw82la6T3t1zJH7SnRg9j3b2XA
pK+in4qEcVVxhfbg6BWnNyb07Wldx/u8JjiAPQzYcSAy/u6sEHvVlVd/Xsa4vEZ0
dR4C9nyaap9xzwTB0c+ownD1ZGPQxm4CcHiF6sVlW69f02hhXsqHqgZKbU11ad+Q
UuelvF2Yifoco5ffxtAUk+OG8kki3+7V8jkJgRljCLNU5f/b070+P60s14Y+DJJv
o/lFrJ6rrUCVys/+XRpEPCNOO3amZKl+4MaS1yUUh6/I2rqJbQ/aEw5LShiQ8Ype
mICgrfPQj1m1fA+V2Iv2PjHCHeLC6Mr5OWxBywHY6zNaOGTiSn8BRUpwX5vjqigx
H0ZrAE/nMcz4ZD57YH7FFp/5ta9ucesd+R+PbGxBxfcrMch3ZK6GizAEBVnggOaT
no14wy0/Nr7CFr4ZjiIWO5ET5ba9XtJbB0gCRDCOl92m9f2huay3AID7UZlENoHh
2vEj9ICjqJHZaQEV326p+AeJA5xhVcLoqZ2SYE1ErUCnrK+26QrsqkMppG+EV6VN
8pQniiPwUPxTvqgjJq/LCWMV/Ri6ha95kGNwcWqrUE2wyeoBTJmSjXZe7n/qj8qV
Qd/qih7ch197twhfqC5mXrSOto2rYHX+LzsI42rama8sqQUWWKgwMOPlef8wopFM
LzSO/vY44N68m59lSR91bMl+ZwAe9p+v4uzTVq/GWnuxBWARtSBrXOFggc8/UJpM
PhSFpzfR9vI+1dOT1f+151Gzjwe3g3eXoEj+S7KsA8VDHFlA+T3Zb+ehvX5LwJrJ
5QNojMF1HczFYDk05UYBONyJ7trxrc0dxVJGvYTZB4NcN2GYxEyVKb/Gzf/G04OE
FythfJDojJY4zE1iXZar/02EWpQiXPAzYnRp2iPpfhrU0hOxzPEP/tKOrQwrILSB
S/acHLpZo9Jzv4hopWnRxTDV7m3f1Qw9ThacpIt+rfqHw4/z/I+LwnxAK/Cc3gsk
Rvg+K3AbSXyebX3fcF4ZSGNDuIOJH0/p+BmQsqkSFIsod18FSJGUefFESsZ+hGWr
rMfRtnc9AXOzixELJEJajwHR2KqKCWz2IaD5j3tqnl3SC+085CEMSqr4a53skfUD
eTAWIFgpSv45y0Kw388WX55Gz6eqfDxZYmlf8h7STHetn2JC4Uj0nX6FhgHaxDNy
+CYNIgqvPRri43jwGh7HzOinUOmie2U4c22izSb25n8OEjmB/T6ghdvWBF+coBW/
jeFVYAgvdCRZrmCLZ6PuvuJh8oFHGuI3+SHTsFWY46G+yXqajR1Crsw+R8a8rye7
oKIqgo9R0dIDCuLK3nfFTuNVChRyB8lBg6cLc2rEeyh8l8nMZUga62X+jNuGk71Y
nFzj+5tlabcSDLlUheHjg+3Uwgv7WOHj5c9LnOAJF4Wo1wI9ItffhkHf3czMMIdq
zZseT07jmvUMxpQ8AIf+SGJrEVOH0kJKs3RMpBmN7IW4e1shqIAHiMEOSEOIiMqL
teTUbTOhh7DQzTUmTuZHYPK4WP3tUyvPmJry80QWVUV8jrkZdsfz/XkN8DA0h1/l
6PE7unhosj8JnKgclImPSu0zPoYzUN4KcyI5ZFg2hM+3k+bC30aG4ir4RnyWzAvi
7K6/HP5W2dpS9zBbepUmWmDVSsqwxxogOOhEZIfSawqGvFU6sxY6dwvQywL7kdFP
BJhkBN/4yFKM0hj3t4R2cy4zUGSfeGRcmw4bSm+GB24lxI6Dozal04D5eOV3u2Me
T+Eztoyf3JNhoGWW93312skcRDnKZ2xyjGondT1j9T1X0FWZmoKt97wYRPbqDeoC
UikwYGGHO3/GZ/NSRmtnCF+FzmSGzJNzfhlX0rzt/LDV+kytyw9yWiLuiZZo0Jud
GSISvCKS8CeKuMJRRWwZmZzCVF1LpjJFwnD3ZgHSV6N5eNgiuKM5QuoQBa4Vf+XG
ojTTfgPkE8+pdCMqlapHdf8G5PvyAh+OLaFRvkjr1oUjX9NHgEUGEI4MD/sQRaMC
RG5zGUO7KlQoh7OFMRIfmu3cT6eT3e2b76JNFYGPVWLB8vU7z/LVBoQDZVyl9VUu
wAwHRvS1XwWzYIZxjuYF8u+0HvLu5c5RkPAkDTiF6Cp888sVYFotjSgm+9Wyy5xI
z1nnoc4VamD+RzHi1MJEYKYn2mbSbdjpi0oBsH0lwIiE5cTkEy/p8NikO0iFXwE2
2JtWNT/GWj99iC3v0EHX4ED2zeCCicOJE/hCFuu+wEHtPsDWiolfuUyItivEFNSX
5yjLUZZPwUpikMGXd91HbLVg2YvunJ2T2nZiH8Lpg0QA7Uf+HNWJB+o437WiWuDr
uO7NmZHOnuo6b0fMGNOIIw03PhXUhg40ru8zuWgx/FhYMA98d+TI9R4L7rCPfOzf
Vbu/7EHgTqk+v0jukR9JevrgXjx8UM8rcUpLeAY2xnQefyARr8WNuXCPl5gIyzX7
+38U545Gt5kjklFGh2GhR4oUzlJLF3AOD4gW7k1I6FKNFfJhJNSUwMpC7CETn0Ua
uK86J7wHvyHv7izjg5gspXRZF3XJb+zh+twsRb2WKhB/KLLVWYddiXmCtdQcujJi
DQ/GRze9myC7yRsKmbO3sNZGA+Z5yoSOI6z+Rak1WF4Z6b23a/XWUgXpXkVBqLG8
i13uN1pgdi6/NS4lY5IHKlzjJbYdK+ajRG6BTEFmnRJkShNYceD7yt6C0YamJWtl
9vRCRLrKzSEyS5VR46IErxD+//+5MF59bylv4sfOIugKeoOt2NGgXzAxjiaJAJPn
eaWNTxdDm3KN+J5r2ePd28w6bkbwbW7Wm/J2lMsf5dILij1Mxn8hUOqfyBRX0DqO
yyTHxhl/9FbgkYJO5anmdLKPfaJuiEO4VY/YxcM/bHFDftXqwvYExAm4sIIX04Ad
DRZtPtQy8ynbV4dkgtlYxJDYy4tXvkIB2XMNUzm1ZYM+q6GGbTmIYBabG+PQ5z4x
JbpuXQizNB2BTvudyauQa4efutSaj0HaFZAR0BFRBAyAm2BPAKOshQQBb3Uytdq/
2dOixvNxQZ1jbKF3l52K0Wa1wo5kkCcTsxb4JqV2lZ7eHMvR0eOAqkhmDxY+C7u3
GXp6/cFkf9MezNn2Kahr5VZ/lDt6V9+GTD+TLxM/JH2U4Ri+GgRz/vHE23yLnLpg
abW7N1npU8IewtqxCpbD30fz4n25D1K111xyvjzgFWpDS3SdtkeJqWA0sVpSOv5Q
y53NKHpvPiFv8Xnk5hlWeJ9zWD85cLSNRHCWxmOud5W1hqhmDG8z2rDF95seHK3D
Wh0hoYh7sBwu2J6v8c7bDXaQzoGEzzXGUAtL8rTvlTH+2rJISxy9ZoNf8EinQWL+
oLTE6+hyzzKYvnnRQxZ7yTD91ex1GvYthX/E2ODdBFkkCuvXntEgi6rAwdY0pOKd
YDQgNV34WDW8kZC5Mjk11ncRLyJe6PglCrIvGnpPm0YkWZvutigvqLKEh4/tJaro
6htnGgum8vWw7u0Gz5yJKYmmVxWObs5nPCmJJjtRzS55Vl9NYfsZ0RtPKM1oXarY
nq6sg6mOS7QU51IQY0sJSYLO3bYRXw3NttqwL2uQS2NejyYxcAcfMyGZNGoqWoP1
iOG1qyagtzReFGJzsPzqoaq+QWP+JN+TvnAyyvLwo7BtEhod5HlbYiuOCcuy9bh7
HH4fGNdtd1oMg4DXrQXZp0laUFRaBgRX+9rU3Re5wQnY7Cl3PlAmXpztuVWmeFLu
jYOmwhMglgQcgbphbSH1DFmSMsgP5syp1/9j6mkP+mXOnRXEnNDRGYGvdXm0U99Y
nyiZZTrclmfIKeUtpIs9knSmBPCyRD1uYGqXA5YIOaEp44p+XFxIu3jUgl5ce7ST
cZ7QWiVpdwc1+av861vB7an+TBjubr6kj6uNjcGcZnX9D3MDZzR6bPR32hBZ3DxG
DkKuL5qfoG1QF93JFcIZhE193X57jl7UTiWsMCjo55gacud4sU8ruK4ENZokdBh6
RrDXQarvOvBNrwyhD6oJlsqFpoHXF0MsdQDLfNMwPdQC9WCaBlGf2CMhmkMU+EOr
V11abhCHzr859d0LPqkla4Dxaw1SBW8GPzNLIku1yHuJ3HlhlI9JlMyspVwHvE36
U2ILODNQMCBTaY0YOHsUi4HLJRpR1BJxjxVYpWA4ByEMyA+RvXII46+1/yt9Q3Ec
Y4o/gsGyQ/XikEf2lz+Z63mgKxfxIpnNgNJSo5xJCFn/CJPaVP/7/1x/qOQ2GvMX
v0cj4ZwM3x7Uj4Aif4ELnqdiy7KYswn8J/gY083kWCDuQM6ZwtUHdxIDWupQ874f
JpXGePX+xK8y4IizUBxl4gdI6qQePHuiX1l92NQ8U2hXJ6gBWemQHGZslyS8pHSs
FmosG3oqiO1ctexuHmWd9JNhT8lhXLEXAFZUCuh2BSOaMvQfcipahWLb6+L9DyVc
nG3e8HfrQAiP/BnyK3D2K+mPpMeOtpY+W8N13eKlovP+JQVIPkjOMwsciOYqmPk6
Tvx+eF9TWinEaQBupiAIJ0mmPJpMvsFCY8kZqKxgXrebfZPbG2ibLLsRydmUIbcq
fieltV3dharFx6K3whjYTuWnUB+1pY0K2gFG0XFY2rOaVV+dKS0yoXxRZnQ4gN6v
bnNJoMdQbWk6yqQr2xPB4/YCdsxdXm0gm/Q8vgw3tKkvs/3CSLrOvxmcDxdCia5L
1Xh4y6uz3jFtQvL5LPxkQlbXba9Undbh4aJJj4SmtiPB007WmSEMKKCgFlgnZ2bZ
rEqbrQb9Xj8zzAaJpu5jmkTStfK+/1DsIb/pXx5Jf5SqkQXKwJq5GUvHr6IB4j3Q
XBTR+vpa1Dm1r7W7JD2JlA43cxweqnvBjGLOMnUIYafJoTktg4k5w04rwRw3eTbb
/wb1F3oJkcC+2uzzsqptyzMjj5hNV6ikI3nwL0hur87VMSjIStfJHmvHBFqMKzM1
XTcjNmW/QyMQHI4hM0Echdpg0xUaQ1fjkNRzDHM5go2t24+ZgFgITqeh8UWTiyKT
J7U05pT1TE8IICc5MZsGcT2gcGgTAgIlWdv2wIIuaqBoOZ9EuVBkIEuOfm4l1dHu
VBG9NEnxamQiIAgrKFfsSG60QssYw+fjoVhr6IWFFhuKEW/1YUczrPpCxyOVD8l6
BBjlQRjXJZsxWJLrd65GtJ7gsWCLS6CYFINN2By21uHvsvw7q0TmVHKGC8aZYcoX
3tqUleEe4DScUJd/eXS8QrBcCsyNbB2+arcLvaNESBSY80lZmukIyZD6llx3kX0t
muNtZ9Oj1iyMyEZZf0PJgSVSbvkZD5U2dLh57GYdbWlD63QpOEdITNm4syPWB5g7
RUOWshiz8LDwtHZKJvo0wIfu2raU2/pw9l1I0RZSXpCNwthpRBvRkPYDJ6Evj3+5
v5rKLc1Fuvp+hgtHmNQQudcVPqwnW3Hkjjsq6SRx/lqW4REV1Ve0pOmKIFxnbBBT
/JaGs+/UG02N4+kvuIEzv2GD1GUrgJmZCp7zt/a+FLKAKervr+x3saVORXGCKrEe
VIrXtayJkdYYUJJ+6jt+26PwRGzN3TwgGpol2p0w8sBjzX9TUWh4PlAPeYdIjYYa
E6aRQ6+jzGKd2Ze8gYUixxWed95QSBz7TC0yPUWHqU1RefAdOG3zd8W2uoBSu+24
VNx0ZgaQwtjGUgIOvaCQ8IugvDTEdDwfffc4GOYoecuHL8B/+1DREd1yr8nozcs5
YNk7B3kER39CE9FsbWhoJgaZR5VIJjmuxb79sP/KeR1yzYTYBKHnUIALb6r4hPho
VpjJN8Pe8SYUMzC8Cshr1uQrgOPmHnW1NxNAjoEubjB+H07EEAR0oj8NRH//d+19
CnRWco4+s6S2Hkr+l8l3NeoIBTO196+/1q9y7AOJUlugzMhg8L2AHjjOWm89vq9q
Whwl2gsjhpIFtgKu4bWPP85rc7WbqXM1FB+Ut1mimVg6ntix2wIDj6JfMOekrSG4
E3j09PYPe3bbieNdvHKLybu5ETrvbKaGF4MMSmmPYsli7uO3LvIsrybeLnt0jOYJ
SNGqs7YqgPtGhd15NHhp0CPUrayiL9oTa18iniZsRfjUm7JtD+PFr9y51146cH9H
G8J7m01wu3AJnSECm1nesKBhi35UbJBAOarPt7KiUGcLsJrXYU8H/Lkpyavs55L3
ohNF/pgvAOxDPGLVpy2VrqIQOd8yx/PBAmRk+8nQPITCdbzcvfVsKoBYGuxasPEL
YzPLYR/ivCNNt9bEOJYSbvDxUXawJZSlbdkr2wcOOXcsP252nrVFpCub0LMijQwH
G8Zj0jH+3krVD6VqnrrRUeDqmnlo7GjkxV4KFrvZkq7ZvS50/w3r4S3+S0PEFH30
G+9nhF/vHkYCTvPmBj2Eyu3lxoqPXfTjASX1qsWQeHsnbiAxbH4S5a3eR/f41ccj
LDe0uB+nktZjz2jtZXt62hO08DfzrBag2kSxUGxJyp8lpjX2dgMLn+2yWI2juOHm
kOnNZ66xfDHWxshctNGS4uQliPNvvJVVIDEq15FHOLkwuBsUHbeH+Xs2mtlRDJgx
0Uji591e4FOu37fCJiJYBjJFJV0R7hMuLVkdzjgiNox6CCRof/2R58OsdnMHRhQm
ZcKKynJ/mazKFUUrM9PKGRjsfziXD5kyXGSToTMTVZH4/Ykx7s6YCkywYfI1xE99
2DBfHfi1P+ao23OTle4pXpebj/YNB5GsEfvma2Aj6NZbwJiNITIpU4ipc+J4Lt7M
x51WBYcjL8OivfbHtfnq1Lt4wDYW5CyT2TLhuvoGFhRl826qg8FbcozapZ/vA5gG
8DhUa6OYvxo7k7c+0Vl1eJfn+Xwtx0WqCNIseLntceKHfNyv4wN1qpJRYUq7AZ2D
rqtP/HmIWnvOCWS5PSgNJX+ek3sbcEiT/pZSpBuW8EmpfRP/2dVc1HCMY8rVZAIs
QJu+dI1zd4/DoBEojiFVy7UzRp3HV3uid6ZL3lE9W6jgAIbNjbhJEBQRQKl9vxPC
6GrqkqSbySNVImxWEE5nvawkug/QnzfRlFfRblp3qRQPPq6NIABxSInY1M+0QAAk
Xsqt46ya56yi6NT6sqkdQe4jmdveuhT7pQDC6skoxB1VkbNoFhdg5d7p/J7/2wux
ZM8EOBNXmAaqwPR4W1Cng0XROsvGMfa7SDOQWSI9FRk67DkdAT5TA3tmMyeiFJdg
OU92HDikajR874R0LLFKLaey66QCzqXubAHhVwm6EZsiBkQDRoLtPqQnEzESpJ8g
hKHJCcKkL68eQcbg+KlNp2UH0M5PxLNIDVTZMSdfNPU6/fJhW+TC2GbX5vuPBoIg
YeekLC9WzexJDuuM0XvsGuaLCGt8E+rrixMegB8+gc8lNZ27sAxuu3rYiN4MvAWs
lMHAbScj9ol+4pjDo37BmMFfqjz1IeUFu0Fv4Ip9W17TXk7juWQXGYipCwSGi/7h
ObHuF3XQTSFbJpeMhzkAKy+2lIwIbH4h+5ZdOFHYBpZnYjVIZiYJ1EzJVq21nDMZ
hxDtothIfCSBlhGnjgCX6cmDsmR/zLFTClRhk94cMnAmcaYCuCjzBH0qQ7PmAaFc
grOzVS8ahlon7Igh/VbGXhAwvpih/HvwwCaHpCNdk2Hx/TSTfM1neo6G3NhgFXV4
CNG1P8NWVU1IfCDGlaGW9Im+ADwq9SXovWnj6nBbCSkO2iCvtJE5zlhJ0CmCPZP2
fIMbZ4N7WVVCG2xWHxbFpUU4lqqwiCDNE2O5jPSr+mK99lHaCvJErzcie8/c/o0/
vwhbXgahna9YApBH4Y3bVII3oCRPKBatoqjwO5MjJ1szwUnpg+mkY/g4gDGajzAT
idQtr/EbuWGQnmRCrk4WyoWR/ehjx/9723SwIf0SfQXjPt0PJ60GPKQCoK/ZUU/4
vP1cQcVL+Ied3fNKHEZ+0pp596U7PItaY2vx143w+mpRY5/sDxhEikja+oRP8Kof
ZuUN35VKivwlYUZxGg0dd0gZygFrhviT85Fa8gw7pEEF+p2atB9kQBAzde+Xnw48
GhBQ3NdaNSa1tFbIHn/yW/6hgqvAtFHnQk6gPXIVYCOm4b0qXMI02VbvuwViAGra
0XfIy/MKab/BPwOhovaKZQrfeEM1CEG6OJMNKT20ZH2TOlpu/WtNqpkm6s9smheO
xKzySGXKdESv08pkszI1sxINceQ2G8w+FX+THMxfs02JQjvMhTsU0LYkL34kfO4Q
DHgELXi2rkOrQS8NPjZ9MbREX9s618eSw2Ws+5T4SXIWb5IpemTafPTE9THqGpNS
kdNw8kdltFJfFxoruWIJ9Gw+vxswg6CmzSXltKhoj/AjtaoIj5YMW2Pfzt9c5Nbo
hMo3i9a8dPP7NzhQNqEYzUUvHuE5tLQCJpoD18ZkNqA+0CtGqIW+tGjRdDUGXntx
n/2W70RmO/xiVZiuTmPvw8gtUna8HmxA3BL3ZdpwP7lmJEnL/Segc8yHnHfHjJvy
mfDo1NU3yli+4Ac9dNUBDwcaIbjpE3/uL727s/+0PmmCEVqRIRlk7lxRlxMW3joN
H+8SSLkM6DwY2GwQFwZw6TPreu4gJ6MtGQJv2bIcF6KEVZoul3TZ6RMUDSe3L7V6
fWuXWEWpjyKRdxqh0bfLtGHFhoEBqJKc6mU0bCcfmfj6kj4DYUzjzYtnlXlf3WJd
+GVUzVKfUuqUC8a4XDRQ5+F0KcWr00pzR3zpMxLSD4qwGX4Crv6P1Hq92jbwaJcv
q5L8fNkCiAsWHDZa3SERT89Tet9sXAW24RMO6B8NRn0lLtG1NzGU2KPAfKFsm/9Z
4yaqi1jrh+vi5/iMWEa2p02E/d34xi7SlzeW+RM5CB+XqDnXDVhYcZWUNnWDRequ
jnBnDa/UqRKL0Kh39f5OsuCd0frwF+GJ9xH0NoEbb5wBcR43ZqKH2NHf6ZVJegOJ
UAyIgAsdNLy1kJ1R63IycIAM0kMLCoZTfRvF6pGBMtU1U12ZTiFea5sKvvef4nrZ
g/wvJuLlZ3/nTyBOUxJV/6GYTEX2TFOuAi6dKyPw7r8lIq8e3DBArYgy1SGbYGyh
6QzzVa10idcjIa9qV9MHuAApyMB2KKAM8yGGhdUyAhMR0rFRrp+MrIpwsZFb9aIc
zQhG07goAJ7NPNkLy8prbFCPmVdYYNCfNBjPa2uGJoKcFL1QKk6zklq+H832Seb1
ddjUKKzQ+mXrRoBUf8s40ZxjzLycK/IDGXIazB5SGnVqa3QICM0QZYtm8ObfaGj+
edDlkFfacfFk/nzMC6aLQr4zdzkmoQnDLYk741yDN/htXsir2NUjFt8Gxd7WT25y
tyElQgVGyMeNJqDR+LzapW7oW1zRjk+4QA2zK8HrlgG5ZsBp1ymdkqbBuNNmApPD
Adr6LcA/bCHPZSLz51rFXspKBb7M20U9jYKle32V6CxYHyyQ8uj3h6zgWqA878aw
wLQjQV4a7ETJQyesmDNiwbmVJtDAW7AtvMTpPM2JEN8CKPrNDPBjALeEXClOgXyn
Qe4Wp8IcunsQAfT0cSW7T4hbz2Tf8GnHhv+r2OxRT9D67e2EtjChTBDFpZkNODMj
326ssogdpmUZx1ihmFWOqmaBghuKEEV0ihetVk3VFw0RpZltth78RRGAE6oJYZ38
KQbDVo0zp4aXXqiG8wdOj334zwC0jWmwpSq7DFR90ZUtyKxor5YKAwTywHG2Ch1N
CVJSoQSuEzNYMBdHb2gIjmEdVa7JCUZXwYEndA8239qd1aO/3nAFVz7QZ78TD0e6
l+6P5MgEWXIfY0epQai8EXgbweVEWrPJfTmO8RMLvsvV/rdCjaRgF9jXern8Zh1s
N4mO0Ub3MrrlCmoYWBIdHjFAecZXmrkfqEaImCLFKdQtbOvTeLNjjN/9jT3FEcrY
lnqKphbQYbWgG88JEQ97QByVrAkTZQotatEBSZMckSSKF73xD6/vn+0uBqTST6Gw
TeCvvS3CeOU/YXI3xw9A1B9IAph709VXB8KNtUe0pl8RXq6y1aYF9XrDf3ALBbXi
fIrIqfm4j5c0IC7QY7BfXhqjUKc83zHTnFY2ZKDQgWVI9Wo1Ei7wukXs3zxqepzv
uARDQyAoW1faZpxZllg8L0L1tiJNHCbCOeq0Ax+7v8Cl6gchJDiXxy4OrnUzT53B
bfkccAqnClBBg/jd7YKJwK27HT9GnCL/xIlvHbjEN92RATMfPMAJGA9YaAuRVh7Z
2G1s1Zr0rncSUTA9fV8z0Q2hKo0LsohcvAVxidQqJtK4L0mKCgSWYP4XniANe3s8
fbWJm+KZerTQ593VKhZjxfTIQIvcHDp8NJ1fKNW+JZan7VKQGEThPps2DvW6GsD2
weUgnhKv6cWrmK5i4ABUyWE210shEUJ787FvZVd7dCznVJcN1pX0qswEVHOzTJGn
rkxJc0TJq9+KjmkioNw/sznO2Cgo9jrA+hNyis/FuPQBddblkivOvcbnkNiylFIs
BgXs6PLg9nBBQeod/AIxIH3wxO825J/w090r+7GiKIcSpN2rdLKdQVkXHwhaTkER
Av50WS31mzNCO3g2kRWFXLtTK6Lq1lN6B0jO1btTS4e82wG4f77vnmKGPTeO8/R8
pOxChBdiH1iGeW/om1frhKxKg/78Utarru4QvUa40uPJ8OEPjn4wgV8BlPdfHo7q
7U/7LEkRz+iKYQmFiYoD547OUXG0WVSOrln++7yNxALPa0b814GE304kHt+WEyYf
1geNAnJoq+XeYlZnJ64akVdF/Y2fp+o5si3aPbC9eXGtlAjOPJ53erjkMUoJ58ti
pBgQ1UwySMsYDiE7je4iKuaeHym8irTAwgK+4hPvI41zZHa7h6wrEsjDHCWek3Nz
N8YSfV7+LfUYcNUS8iWGbKgrsCFIMtu8X9BbjuEqYE7qCM8gzavrQRUdbht+baGy
ZIz8290qDykEpuijtOS/5LWCyNwzuVpN55HrfFkHIm9N0IA3xiZSe3jc3l5e8DBH
OFbhv7EaW/qiHm372+mgoOReVxN2/NtN4IgUbwAGb8c3sXoRerZfcAVwSpU0JKMZ
FcsYZoKeD0K78gRyZk1q2EREBI0/jCqpYfMzyL8pntMlCp/xu0BQPOnS8hvWO0My
Bgrj09MdTWjcKKS6V/cCvRHoozSewdJpF4LwBDEexJKABceqXK67eO7KML/awVkP
u7xVNQTVfPOeV3k50r+OAADvZLbVfkL2GdQQuvsMKUGyYRy81LFZvmgnz1z/a+6p
ZgEt3S4N29qrMwH6dKv+A8KDPUdHOyKTqp/31Mr0z9Xhpd7ZyGYU3c2K/tLn24q2
pxZkhXNFO/e3/Hyb5T7vrNyG0NP1cgH2R9RBJTOEPnW5VFVZ0kAlHobyK4Uovu9H
+5NO+P/6O0DCgbrgBhKZ/J+dvjYN42R3Jl6S1m1TVhxDxGpLQ0Smfip0e/MUTqD5
euXyMljiv8nGxSPmSZ2jq1mtroHBOLSDx0fizkzVxy83Lx6ac0c8g3+ibOXbSIS1
Knht5qgdQZyOtp+ncqU9qFjefuWJWlteeOZe/fSNLgT/eqG/yc/eNMJjcWIXHbFp
GVXLTfacwlFEDEX517J66viE8ICV8YMgP6voZ1E4+7I+DLSIo/GXm7M0V5e6KEz2
2bIqd5oRCloirjs07lqG+xZBrT/grgt0G0MdD9ZyuIBlC8DECbpMmFNyJGEPPYh0
BAV1w7HYdG7HUalxZGpY8mztvrWSPJRE3QhqZ/lcP8p7Je75NzHaKF1gMF/u9IED
qzm2k+dYc+OyFaLUkjUR3QY2gppWhe4LP/29hkbiKySRLG9csM+Lt3XH+sVByqzk
azguGbMVXefAd0rkSW0fYjKjbg5scaA5UWhq5a13UKCU60E6MehX0ea48kIpQ0l9
WJ3Ntc7nnw9IBL7KILn7k/8hqjQ3hiqLEzrgMCtxJ5KGWujZXy8Vbtd+EJTs8NBo
Gx8adCBpnBwQyb0IxhCa6AwNe1bFxA2T3Rkz/a64ZpC/EEnUfmyRb0KnyYgMSxDM
Mopjr7Ch+E0KalmEKX+6eup9uUp6Q1fQMW5ru332A7oeVnO1aJZT5p1VoCc7NID1
8XS1brlxIDCEFYMUkSF6XlN7CiNLekibJBfJpJvU6RhElxEetzXDeNiPevam9108
jg+eOa8q0y45aeFqsvwac/1k72WhYSKTIxFdEmh9WpxOLpNjY2FRQxSK+0CuYxM7
wpHx4EZ+V97EOxYtxbwis6Orn8JJVJyp8djsZv4ytuIjINUeOnQMRgB7JwTLQQBf
zlT8sXA4CkgZ7FI5Ho9ah9sIjJ7yBgTOQr0w5oNFgs3xFlg8jIrw/2ChQlk6d4Za
HGDY7pbJy6r4udEpStwTAL9R02yKzQeSaHftUeYH2dqd4ayJg9k5ifnvhEP0RW68
FnTXm7ExdMQsLQJXBdInG9XcjhbFUJwY7Lw2Me0hwCa7LoBICZCZVU5mDWp4TwNC
ENDj0ieX+lT4k03WY8PeC4uQC/OhDOYBnHtnh3dzV25uKIUtLCBac4O+soYvrSmB
xl3sICJz5l4yKm6dXnetA2TL56fiqcITHKvO0nQlpcneZEO4M712g9OiVr2Xudd9
SU5xsuOHX+IX4VwI6dN/61PVYc41Gjd6SnT2h0+onD+7ORtS7fnyFkSf40mdT67r
4+dfueqRiZIIbc4mMWfW8W8MnA0Umqx3BUX2Q+sjIspZxKrVyukIz1Nm4BD6ub1H
O9auJXcpz+OJ1qhA38t82NleZ3nF5DEF4VqiE+n9BRwjS60n+8Z/ujtC+wlwY4pi
BZpguRAqmNNomDLTew0m6BLaxjqTldYi90dEgTp7GL1cIlLMJM2/AWxcrwNzTy2b
O/ma6Zt136nqgp40mA5pZi2PBuucP05eYsz0rPv9tNPHa6SGCC2F21jdpcel5zqd
2LOrJ8hHEQcXZRKOCfJJnyZoC6cPJ3J6kjJJsf/v9mfGA9i6rIFMfnCz0G6WBmdv
idOBDGwYNF3KRBa9NQNY3MxWUMoaugOvwZ9gFvHpHge+fz2+tAh30pkbIRZbsKHK
BD4F2LoOw4wnLn94cIppevVMn/EfZQIq53i6xiepWs3QC/CWl4bcvmkkp/8SoM43
GlIUJMP5WXoUxn+8tIBQI+0IvSH7pgbvdsDwhea6wwdaHcR58G16ZZWMNrYwxB9/
pH8aHNeHH1RAYvvsV/V5Pc/6Mnzd3lIdLd7qfW6d0aJpWkZPYkZES+r9uVT/tY2/
Kqn+zTzAv4GOORUzMyn1QvWQ6awsL139ufIS/kqcXBSzNmZceheWT39EzznjZ/6s
JrD28yqoqmmwhKaKprSPUECBjwBw+P6bzCzzLcmzqtCfG/3pihp7HdN4joKJJr3z
zG9AfPre3HB4TMKycQ3VHKiQx9pqZdRc8Igaw0otU8jtVLZ8fbBMmSnoJQ4yFQX7
dfcdlmvHuCp7OmPV2hJYw69eVguNlfXQIXHwqktDmaKN53MoQhHw242mqPlEhTRT
PAE5SZvdo3+bLqZOnUDufy7wI23GA4SZmnWhMehmNUykeJt+nq+z7H33990JkoTh
MzFYjcYAIEe3pI2XruDOsvUXHystET9el2y2/BTjELUxIult6UU6+krhLHui7sdA
6IrDkogqNsVocrFANYMXe3f58d0/JJM35oFufISPhmGs317qCOIFJcj1+J/rlNp6
5Latrlrqy9cKfiUKdT3zwx5lgklxLtTRmIUdbHUa33OjMOs6tb2DSb+0JCXsYIfj
cwAbxLCW6Dd++XxPx2q6/gqJTZj8aAYCuoD3fNJnr3YIVFlVf1Ed5TIhJ8Z1PFQC
C1RT2K9UAJRaeZskSiRkXSORzYG5Nj1PvzwlP4DTtFE8BNyAaA7w+p5/TaPNfI1m
Pwj/GoFSMXPQmceTCbKiIZNFK7bD5Er+lg7BnVdpw+Mk10IRKYwHhPkUhQTVGcDa
V3yq2xycwiCWPeVlGB9m017yNZVQdOrujaab7Zq8wMFhf7o6IwtYTBstF658rod1
ECYPs+x8UkGSTTfPJLa+nPj18ZlroPsN9bSSMA4djQO08LGkZMRMI+zgVEC/LdyD
UuDbJfv3uaYzvdpOqHMKd7fg7LYBTnLLVV+eC+gHBfEXvjk9hEtBV5ZjfpNR+jjl
hWhLV+0VkBUfZpKZ4L4YnbunvQv8c6E9BKyxyPSKJJqaBOxKihxWy9wIaeGH59Re
RiSYonQWwDQNLaH4yfrmG7CprVfh4CtxtfsmIfhq7StPrC6A040JqAft5t6xmad+
XoJ2FDPlIFiA4MKcFTezz61sOBgoI2pEw2+Y2NwXyEI5JOqHOZ+aKmQUp7OFp+5n
M63AARi+KO8ccBjDA9S48E7IFEExLtFti3vJWR1HaY3HsYqEip+MMy/FWW70tPTm
tnRv+pSiqOiSWaskyD3aMkdyKZ6GO7J78/xZ0VNHFHh5yEY/6npBqWV0fKlnX0JL
ootgHZ0gB54UBS4OJbRRt1D5pzYYUaAUVbdze9w5Vykh8OfhwTfDeJnhmG7MCFCj
3zD/jOjqbw4ljnQnlygxNUNKQ2MEXgkZb9B8YYayEGPUCA82v87P7DR5qEzRi3rz
u2zj8rXxZ3M0g+WIP+kN55d4Yl2sgi3bCUH6sxRZKVhfIJ1uJSTOO5xX5ArMnrvV
KqAmoPwRYruAsaeQ4+n7LAhjP+qdkhEKMHVzn+zBUEAebpRVWLJI33y9m78KXHLm
dxsbv/TWg/2l/ZYf/PSSfoxF/sui53zqcIjx5I9BbdxMepWFmnTTxVZnvwGaNNNA
8oeqZRdNfQFdss1GvMdtmRm0Xd/uKKLHkWzINPxeFJp1/uiEtlJhHBmJEGrG+HDs
eqkX1HSE4TNMmJIU8cU5FdQn9ueJkcpght54J1xwmeodaO/zhl271ZYovPpVLija
bZ8P36tUd5+PHOdu6iT9CcnhD/chzy8xlTxtfIHPLL9HIiOjHXnUbZ60E0/9gpVd
o9E6+x7VyuhWzyBCUF4HIOqMh5iswetJKf7z3GFrZUDtPw/W3rKDo0bwJXWN59rU
UdFnzowSqGJ4SfNycyvesPGJKkJ0WcaZW9glkmPWZFw9IwSA/Sk9erOwhcmEIRWO
rOtPevAcuyodWplcUbAGiDivkkBzzFoN2+x4LRYA5L4Q7hp0AZiND0RrukRV2lcb
MPhlAjQEd8zIuZ4/iTHdXbSlJ8VqecsdNnNb/Nj2JYNydE3GQZWtN+5kK3t7HmhO
9Blt8oJ0Bc2iyfauUCrOxYNmuDnz60gd52hoNNZqsnMlUyQkLZopd39rA6LkS0WG
9M2QFZgYSv/7AZYmULGrDU8DrlFMk8R9Tz2emH8acSJjdplf14y69qK0fxoFFDhX
TbG7cOUMT73DeKEgi/0bpdhPw4JeM5kx37N6IjuDiNl9qgM7mNqUvC2tG02ruf5y
EN8pYMbBqIWNwBfS9uDzuhj9cTCy5NpL14jsDuQnEVcjICfyBUzM76IYQILkt4lH
pud2cimPbBvQtKJNdBK4dJ+J0MPDzZazQY6x64TTIDz+FgZDvE7LtjT0B5wciWzL
oa7ZHF7yqKFPW4aPqNL0nqLZhqm6DsQIekiXomaclW6m6HCGcB7Vwov6ouhBh8yr
pHHcroAGYswu2vBH/Z4nt6oByVabikPkNdrHNnmGrI5XcITeGaAhccQx9XIhsnSY
EutPDNbrdoTi9AV+4JqcpW6vCr0453LaFbq0B0vI5TylHNG5d+i9IETaV32v7AMX
a+E/YkWmSPdgoN1PcG4cd5IGGLATNEHnql63SrVwUqR+QN/o3YIk3LyU1Go+3qEm
4SjxHb+l1kLjnARc03gqyOg48XSkIeIrChWkzyHJOm/ckm+JfOReDhdGX7Vi3KD9
eDcYGGmXT5gPQ3oeP0TB6ussWJJePoOgY1hH2HsmVIn5Eu68z9EIJDb6uo/8/6X7
YXE6D+CZ57+mardNmsCDLTPuSxVlwDZwzZtE9hDgR8tMuhc5z3IQ6B1hrfNbHPtV
ibEMgg3plpVE/grRgn6uyPPBM/hAHWoQFpcLJEtT9EBnGuxDZGD102ZaGQDPjPVP
BY88aFAJr1JXV6bw/M/s0wWh/9+RA+maCE4JT/HUUMSQc9EideXd47RRKYnf/zXV
SB52hNca5FEyR6tJ1x6zzbkN/FCLsFQHbRnU3j4LWV3o/3sKBDWkRzVWxclcjc3H
90ujReem8tm09UFuJGRSA7sLzNC1jUjK83qCO2gBuFwNcvryFZecLe222PWJjgsC
MCGZOLZF0lPwZHy9jHbTKwLrvo6JKPMZjtKepN80NYYGe9nd0JC/VLkxV/SZEeyq
nBFLZTZUu2+NF8AgjvL636+GKMc2IUkZrAwmCAKR+LaVeawDjF31EBogmn1/wKMu
6wCZXHHvbkv6qnZQf7jWTYXezY4NFtjAMvspMcQr4AnKnX/pyKt8NxtzTHYNfsn2
sMxLyBbQB286RmhpNXRed+L5N6U6TkjoXLpDSxNTbxb0Y+AQeNITlXkj/pzyfWZd
3GmPzoC1nmlS3ZH1JYDLGxKQpbm1b3MHFPptVzmP0SyMgPT6WDOAJYFZ0SM3koz/
I93mMGz2bB0eNX3YGkA4Mm0OEVtE061Bk7HuwiEGuw6BUVoCnPvzfEoFH6JfRb2+
neBbTnPkjvoFIMGz3BAGJ9ALTFfY3PXHXaT2w7psK9kcu/iTIWXTPmmgl5fjRpJm
+P/sO0RsM41VE36vELbv5jomo7TrXCNV+E84um//gD07yf6k0wlIFQMUVyinXOD7
bMPQnKL7ni3SuoitI7RCZeoXLH06EzioFn1LiFIuqIXu/zyFNVn6bZdKPx5ARH3O
zqit2C1PYma/Ugke+F2rba+r74QNZ8dJLQM2bQFW5cABqGpJBxLeRzgNsH8GWc5i
lMdQRUb2XNV7Vd34bPBRHGimzTgY2dlksKIAk7Ge7kymTN/Y7w7YvmbeqoZWlCi8
D1A/HrPsrVMhm4GcC1rDZDDhxihbk5kdFucYFqMFs0OysKBtzUCRoK1YB4m95+E/
rkrqLW2kpYj0bh+FFVNUYBTIWKiLRzQAG6IDhHNz3bCPSvUe0CZXwxr433DhgXHd
kVmFk/BOXRfAaRRE3emwpTtRHA61J3qUx7YeHrPKN+7LIderSI6dWbXwsKLzJEPB
ACqhNSjgEFmj516kjG9pjBlKvHk8fkPNH7HVk0h+vlgnzeu3wUnECqtr0+bDurG6
RE/PowNUszVGd4T9Zg22OuN9CaqXHjeyiiqu1zS+2t5cjvuuv6mosgd5CPUZb2uh
aDflYUwn5oyaL5ueqDMlsngSaq95Wuzh1eGvKWazaOMsOZ50ngDcFGnYwYa5jbJ2
PZDxhClL7jpJj7/1xfHniJVhYbBgyvNvqSNz/IrhccuDAjK1EkIZ07E5bxI6rRkJ
TSG/+dtaspSw3TYjNvptEie1tv5aGuskT1aXWIOmNKeqM1svRkLaG30habzzfwHA
2czi6kUulD35o2+8HU432ggeVhtaJsDBZGb2ckTbubB2JUmIZQRqYVfc3B/qL/Ge
gjXffxrKLNM3CxiBgJdOqcXNJfMaPY4x2fC0w+DQD/x5pWUWRiz0F4MsFTLPOvUb
YXYn/GhK/v2p8NZev8Ngnuez4WC+H7w2mggcYoN1Ef4H+zmp6sNUPQA9DG6X0MGv
kAg5vNS6+88QkNx7Niq1obg9omEqWZSFjXp1PYswuX5V0OjG6FJiC61Ss+2hSsjk
R8FqUDBg1YBUDmU+u2dfBETOlbrZKrsxf/6+nzhObA4Rf82aHzXNK1s2WWHu2UIA
QdWUFXN9sy98VqW1NgAoVZ+EGRc9Zb0iwqlaLAa4Uv1wgEJG+Rx04RIdWengD9RN
nSwc41B1MqeZupiAFOM8WtnLvmuKLheO5VwBYQ8/rPTbXtwEGnGtMol40nZHYHth
CN14MX/nP/ec14gpbiDMZpvVpeLSPupQg6N7m1dSPJulVhG4/WME896/O6FQ1hxm
mCLYf/Ptp4AnZfZKb9eNtHUQQDXIauxLh3ITGGPIxaE00RYGnT8OlIf3SUlglVYR
6lvOqGN+8TZgDi7BMu+o8sZtQ0oPaP+4sXyx8LslCQ3Fk8T7+Uj1YNdYD2mOp6C+
7dKthUCWNP0ZIPOVlU6eH9D6efulWVqr1Y0Pg7rH0Y09IguRPypVrac/3z97KdGB
289yUWHP+axXg/2HIrZY5VPrErTPyJVLUirdhoZbUC5V2uF0FtmSWREu+qSwp42w
q9yw9iSQ3/SlhSV4XwqAteA1U8/afm28HAYQg8GVQubznIKFBX2b6OeLHOhDEkub
T/brV4EuJaQfH3sCcJdw51FpkF4WE8LCiYUs06x7il8Vg1FvT7xuSCPlEv2PYLHB
uJxp9BDOS3iZ7L040+GXTFo0RqEfIhtI7hntnwK0213/KPXyMN2L0QntyMOEW7vx
6gHWPvEWaFsdvIkfQGZeKCJizRwZV2RGFWOlQr5V7EY57mfvYYgWUkFOkoLa7HA0
AxpE+KU3qc3UUZgesW5XYsg4DqfsgNmVkcGE7/pCtlPGjmVo7pZsUq1ZPCR8GgMk
evq0KKf4bEtr305f3h7obDUDIvVDCAIBou7WxAqZgO6bkv+kDzlNdEIjM2Un7hb5
vdgnxi/IuKalb7yqFg+GjzpmoMo62ddQNSEcBc0Ds2SkTBohQIKo2WKlxKgX8lxU
6my753HY6ova7GUyO7leHrLI0dCCRjNGcNmIeHIvVdxy13qk1JUSgJv7F1Pp7HVU
odVV+ZvjG1MNSUwWY8zhYwK6I5nSpqIziInUCaq2QYDqjpEgv/Viw9LvFGSi9nvp
q4sPKP3rSHZosTnRxHBdgORYlVTIdp463GsG3nQxIrNs0A5if4mFq+EGDFgoNB9o
nV+yx343390qpeCKQpCOUV59liUzdVUV9UXLs6oJ+5IHbc+12DE60RrP2bLV4Iy6
6Rl3fWhQ2TzlfuEGDYUMrlVjxhEN/+hjLMMKI6CLz+Ht5KznuGtfR3DiQIliAcp9
EDBOIvI+Xgy/W/1z0jf5qzv0Uyw9qcqH7T8R38qfsBxY1YwfwdB6rKo7+c84IXo5
LpW4lJG71JGlNvKHMXaZklqXdsCWE/12IHEJNOkYCxM0IUfTxMJRprsRZd68lEZj
XSKpkNiCoDox3aLpAyn84w2VsHwG776f+vn7Y/ZdXjUMXmK+u3xittlSJCqlwD99
Ge6W0Mc5EO17WrO8mTrZpjogJVBxWvuqNRaCP7ws6tM1lyoSE0tVScukYBL1cgGR
DU8hZg5B3NQfYq/gOqM+6SaLNizb4MQAvEjfctKafdlhGHE3T+NkM6wpGIUq1kYL
M3pg8Sf9GjK7TrYrs5lJp8K6KJNDiXi6jc6rdKq9I7TXK/HplgGP+2A2SpSxBLzF
WhnBDBWMrCPwyahIRJICXWlYZoVr6ovl+62Oq9RhV6xrxjDyqwP4H18KUpm6FqDw
m84mfXFr3p/lDO9wWqEYw9O8zo+Amui+9QtxQINUyA11TjErGk33TjFbxhA0g3dx
/eQAe8NRbX1bm9uTYEM3qVuTn0ZOAGRnmjN4218ViU8oRt7/BbGFC9bnkjnUIWoS
nRwYmGskCaZoNam8txdtQj2ry5AYmNoXsxmKuDaQsPCKoQnN/5FmT9hBJdXYLOdO
u0fZLAiuedC/6As8mFiihfa4SiceAmE6CQ6ABp8x4j+mv5Uc2gMmw2FtGP4Os8uk
kH20HV010+PZxkzHZP1fPPixrwuv1l6qVNs24n3ULCXxiF2ARxwn9hS2ou4sAWtm
Ua+4GxD61WV3fZI5Ka5bz4FzxAGrYTvRx1AgHAINo/xCX7ocfhAC9hig65TeZzkU
eHGeMgDlnPKNx3YY8594T0xWFzqHmZzktzWobI6l1jZ6csd0A5uIrMWkVD4FteJK
+GgZuatubqiiOxXR4iRov4OK5sYHezCazsM68exeu3pRdE7mD4MihqaERVJ1TALm
uv1BIr1864Gddw4bJlGOua6bpArJx9aJgh7TaPhkIoX7b560uMHdXxLEz+CfxkFE
23iKWA+74rjmn3b7IyjJXEMXiFYqSLS3m0RFRFv2LnD2KTLuPn4byL7A1C8C0ZSC
qsdWW5UtlJtKMglC+govqq6LvKHRH1U/CsDI6HXZpFoL6rTL/CETxLkH7u6irIAP
Mb2jPq2NiQ88+avy0G+DUzJJgOLmy+Q3Yn2dZUVkXVid6KZQ7qPv5ca2taDVGIh6
xpxLmkn4+9p0oNqrvd/fskdLEuCJtsh3pS6mbhTVPFNf5aZSyiyOxjV7xxzi+VP/
EeiiciUMDxvHkDmo1GGLgUG7ytJaHArTKLTBu1nhK0Z4qTTbTDyi+fdGjy4sWc8m
Vhg4hLNj0cx58qF0amCkbVC6Yu2CQyd1QWeSKoGPC3d244NSyjt7rXhKx7ynVjzE
/JvoEfu2VrKZIRpV2tWlWPfDgrTWqqvLIe1aZMOofx1f9RrVD6Nwqu6YVswSci5l
KTj6HGpu47ir2jX/p59aVDDmmWJSjGWeql+O6SjMmrOc4bqBw9lTvb1i2qJeARYu
V5l5TA9apwQIKeBKQQWmFhgPJ+GmdnTWztPYHlt0nx0b+NbzA1vIvZFp11PfTUOk
O2Sjt8uLE1yOPweHHvKGG1lpXyw2SKklgsV+iENf5YooAALh1mzGOcrp/K/cGgeL
vU29cKv+b/oDz8cB8bfNsjTG84+TSh1Ns4kd59T6JxnrsUHKqJUhP85hMWvxfHO0
UrbY9xHrwsItrboxlBgR7kKr25BQdRTR1I5zpmmZXndK+UA38Hxf7/kscLgUrgqN
F0aQWUlchPzvHI3CyoTWF5yUnJZT9ZrsOZ3Z1KzOf6JBhoh5WrhWsnf2weNAwwdD
RdiCxgWdNqrAiijQFff2RfNqN4PXwWfxjYmVULC7J6aNgQau0or7Vif+AVoklOtB
HgNk9NgHcSYbpeF3m8/8sxwBlDvB2FS2XKMjUTYTKTUWg5vUBOF2UAVltM0e/NyC
Nrv1GzoS/C9xbM7yBtW/jebUvd/fPtsOwFDtkj0beTS05s0Fv7x2OCzSOHONIaKf
i96CHR6R8udj26TyAE8/AhYW32MsgX2jpM3/BsFvS+NMaHQbM342TSXvXXqbgPZ8
OtwNpTJFUU5GXtn1O9dH6ltfIHF+zerRratsQPbnGe2jITNFMzIh9DqAHu2ANDnP
FeFAR/8ZvAOznQfo9ywcxjjvAxKoi/Vc8S2aLO8vDwxxiFWNp07dn5HDFQtbThQQ
df75cjA2iJx2aXEliaTY/yLLZQJ0PQIvzF4QHw5XitbQD3bu9phQYMve+z4R0XDv
vGG9232J+7b+5m+iHfivZ7pgLTfxe6K6zPZxsacLGGAU2DKmFhPldgTOtjztVJto
mdndaGQ/VkKa4U8TrUNg9JwwtVWsSF+Q6uNRZ58CYrdpl+IiFQTANSZ92uL1Eadi
/7cNlplaW0NJm/uxgn7DKTg/hhjCl36Q/1FKNzDFhXNROBPMNcNw8/EY+MAj9xqd
8FfJ6xBAj5crmfLOPSlw35jvoQe79XtmScXVhrSaPBJymnvQG+rUIIYss9fLIFQ+
dqJQfStyWp8aohX1FBMzkLmRZ6wD91uweEdKw9UMYygh4FnuaZJYn4aht7LHBKO/
DcudWwpiDO+JL+/IlT5D53lvZN1462xaAJmVy+m2DdpDTRzGeGXLCV1VQGsB6+lB
9HBYoXCXD8JDKSWl9bC1W0QEMqCe2DuT5o0Ucu7zPXW2GLOlnwzHAisSwbBpMdal
DzLTrnUYylaNXTaIrfF46bs5pgby5bTVuB6NXBbJ0pRvL2H6aQ2D2n+ry3YWi/SW
VAhQWPtC80TEEPE5o/z2pV/c6BMgMyJ0Zfy85SX8/rphABTm6URQ8emJvsXMdJrs
oMB5IKANkqJSO1FoYC788D7Jmi19aL20Gk3daxg2yOFVC/Y536ahFAHXfovSmdPh
qsmDxSnx5SzRUIqYyUJiRdK5psUGv9mvP/bUzEegBWxsOvMVqW9EBM4Sx6Y0DfFB
KhOTsrYWwliN+bbwfykfNn/JTyNcodvvc2xOp7atnJ+7DewywwJMmzsZa7Gy7jTS
RFwRYIYcvr89JPyjByGACZrg9djXsJMSuhCNBsPK8fozWnD48PFZJgG3ZxlmuYI0
kVLZE84jS/KtjtGYREfit0/+Hi+JVcF2PaKjVGQ4jzmsNFJYcq+EqhsJvj7OFlUG
8peQ3Lr04f/kX0KwRVW1DeISanWe7Eaab0qdb5H4OZdUxePTWCfPfTXUcn4YX1Ig
tHUFia5OvK98G5gi75tU8/t/v6YQqfPPT+ZcP7Cn3K8Hl8l5XGDC5N5F4DPyhiP6
h208yFhraFriikeqNvcxv1FbzrWC/9P2d6IgLmZGd4uCxu0VluBZlboIKiSgMi8Q
v6uh2rnOJntf/nzGEMpDoUxVv2F7pJCwpZzA0HXqc2Ey4Dwxn4rw7tmXm+kUEkr6
1mzc9YXDC0/d/1OqZHlSQwcKz4/ZvI6rrWPL0aqf/oXoqlfQ47VaDh4GkbUcVnbs
aNAhO+BldoE63MWX+zCLUA+/XUUQOOOzfzdDyG3LPpFWNhwbpkdxr415S0Wr7ZxC
jpxoo9WSoo7Mb3gPsvZOg8Uqa7A0EnOBdngYVP7lc5NT37rKaPx4US6/2lDyvRQ0
GYhVgbdsd7QK9RCxUTIYaqdil6ZeAADfl/T8rtJIM7MI0oETrsbTIyOXo/HQbsH+
CetwvCTkA0F9cn5CqR5ak/Mg7Pyb6rRbDBxoA1Y9HJWnpovAK/r1tZGT9slgBXDI
o6lRC/keVcEn4TT/XwmACz9XwgfxtB8BfLT+IxrPJA/xRzfBgdvuva/WTh8vRUgY
06xpk/aUoz8s6G7/AtaJkdXD89bRpPSl0qwkK95qTrPSLLkHBgozNLGH+0wgwX4Q
OgBNZTySb1jq/YbX9Yb6tPKzrfsuOwj8gimfwQU5sSJfe8ua9gwlxRWGGUFmEpY4
KYRYdFixIc9xIlnvpIivPnJisFEm8hSZipIvwdptXH7xjOK9/P1qHMIc+b3WmDJI
0GBgK2cL2mDKlfE09KdSU7MKO3p45rQ/6FTL9JNGlt7tmBGn2oGhYuDtAmSWFkzn
U0FOeZ5AEU1LbMGY56+puHil6ySYZwc98reAgj9la8r+Q2YL1yqxqWui/6cUCD7L
6BQrXWYPz9pr/knAclKcr5m0+IiqoC4ln/s6gLXGKaZZkkY1mTmFnCQnB4ZTKiA1
UPAWaJGYLBYPDJ4kNXd4GUW9g1lKJUtsEIb1/ofFaat9mtOWuaemHmTc8dq1UmGe
J/qLXY+WMmyDTvL/KSMdhte8PnblLQ67LPFxjimZmekSzVx1/OzCQ65+wWbV9DIG
q7lTZ/bFbktYhkGK213OoNtdBRnoIU+v6LTKpgHBlAoKGqvXiU57yF0xBpNZGbrV
k4vPh1Xrh+WL1SHpQjzo/SA6jlHew3bq2thyKQkisbe1AmE3ttpk4ecpNlIoE+pW
qGxQji9d4ac++/1qktxqlmFqjY7FwruZG6MqdCRT16ZS1V6mfw51mQ9iGhNJNbDO
t5ImS7rG9CO0qw5/axiy4eOjqwDmEJcKosQgt1t5m4OgUrn2Sp4+CLlnLoPTwqkJ
h6leDoRD+/+Zy/GtcI4fZUVcAPAE5aCLpL/hm2oekbMrbCXDFYIC/RvrGXkor4yL
6rEGYGZMUWCjung7NTEvohH+O7FsIxf2gYgek9nvXcZ+T0kSIn9hMcIOsr+NSweo
NXfQKZ7aVz+3TTUtbjbxpDrpu9wjDVOOosEss+cOxwEBu5uYkdIYlVpO1qtjASnK
8NZclhWb8yoEemwYG/aa0Cj1YizFAvUWBQU46cF4iafJwzS5/ZceiHTyjnF8Ilta
40PzjBpEKtJbYerGyLXcFbsYisWujzIF0Zvw8Qf7txhWRbVIHbG8VoX1fzoNEA0R
J6AouIVxj6ltDe+JEfd0PiC6OJIUOyXoyfd4uE+0vILkBoJTnaPrQ1nNcgZKXFL6
u0lgcZgzc9jATfHWzq2zVoCI8kunziXDLZuPtIZ/61JDEtXc2bvjeebMB+NmYZy/
N+wi7G+6BkX5dBvXXsVFvAjP3d2EHqkMIxygA4WeLm6YrFY9W05/p6etDnXpszty
r8ZuiGJ53Vk/lsXHAzhLhIPSlC8drTtTpgCgqeG/i42gUmjo3/0ERhadJvfCk2mU
eQuEqk6erwRtdMpRbLT4V0tM4/PyYkXUk/O6PQSmNydSyMIRo51+gwQre432biOO
eTJxHipz0LFe9TGvbh/5oYxIrQuFx3qXhUO4V48mKiHWzmmokK+pN73kUM3SXlTS
Ahemb90lh1w1Di8zM9szBcNGRi0r34FyVSv+OKaDsu/gYo9M0prGSZhMgV3xhN/9
n6INFjbea4eR9piddXmCBJfy/G8gJr7/TFLLWGYSHZR8zKwmliGQj/2JWnvCEONe
5Zc4U1KnNYAy47YjkZqe9TP5ujmf6vb8e8l21622LmnhR31YIRSm5bE/59hIhfle
58av2vaLs2UVaCNDLl5oes0pk5wEZ8zySvrU4uuwjkKZm4/DS/36GhVXr75jKCcj
6lkJDOpEUdkxPQUMtnbbZAk3oFxH21cWftKem/RlQAXVfoivSRtwPWdr0ibtF8wg
+XMVsPQeQ9/W38jjjHELkV0EVU/Z6hNYxRjUo/YVcUFWxMH/fMNwdbXjIkMTxihU
t5+75TdrGbGUEZiLCbiHjIfsM1m+eH8Fy6YJbdpRmhvRSeu7UVW0DpgiDYhKJSRW
bvZ4LnndvY7OEAnTR7sG4zmSUC+++U71RSlk/LPUMozabuGVHWNvbgHEBVq8XOqC
kVx/yMpqP2xgF8211cRELiHaV5YKDv8J8QIyGVJnygKIbgYstrh7clGoIMdCld1t
SLQMoqfGr4k6IwtJmsintGupB1WGWBt8+9qlvRcUMOpEx2Fwm8QEiydgAbwHZuij
CpRjCMDY0vsPlZfz6WfVYjZfpRG9VfzKu+INlSiu/BYb1TEybc6AmqfJkZX8dVH6
OHBnf1OKN+mhGaHjsXrGv2Nkz4/+ybgKINjOY6Wt4dZmSWjge8FoVfSoGcoAEfXW
2lTou+uCxMUN4ZJeYRyAQVXaUhn9wjtQ4ahPdHv4sMyKWegWb4nNEcB1dO9YbQkb
BkOAT5pPPcSdqXYiX9IhdCIDMlJpmMeDch/GfeD02zTNCNZyFGSApQJcsKYayS3n
CuFE+r/mYq34oxdZ/1OQJ6z8flg9s04Xyg67u8lpCVNp7OkK6PpOXw1WQbHDglfV
U6qBT4Dd0cObIYN6tBXJQQpsax5v9kjBWZCI/wgPbns4DPLsw09CIj4WhUCZHk5j
00QlD2Juah9Qzl+9vXiJQ/pW004r/lljbuhk04e0gj4dZLebiDpUWHnmF0bkc+fp
hfMd3TG+Xx3+CZxVl8McgxsUAENQhdhNh0uVQGk1Pg2Xg31W9ExstMmozj3Tvxwa
gfOjbgMdzMJKc7AcdX/g2Puw2+dC60k9+k5dtcyZc+jX0BMvsTq2My3gzzevmHiM
zltx+l6fxvwmzxfavv8UOsQt3/q6BA8SKj+DFHllc5MZkcrJdKAXDULAwkmteOoQ
t2JTA7b7z6EbiX2exZW/Aczc9RasNsLgWKey8iry8XStQMZOEVaA2uKrDggQjjR0
yIWPHIfOHQVeruZceJBhfK5KBcerLBhHRIxinTXyh/Oasru/AXmPNf/wRG0OGHgT
PJR8uPUlmJo8Lo7APj/Fr8M90xYDBK2j3wemTrN1l4ZinphHG4pdF3kPqClFsYbQ
MpZCc+fu4+mwzSmChXiWcJ5BJ+ey2HzYVk0L5npBBa5CUBPVXIyFh1mpJuEHnvPd
LI6eMj4EwhpSy1qVRiNPBwXvA/MP0VYZ1HxPCu2gZaBOAqohBsvvxcazkP6D/Hjn
cPvaoIxksKPhk6v+EUuvr/eO++0bF038BpTbo1i4yp7ZFPaFXmbk8NuzKGEEGVj0
1HL56YdyWxDJkYXtlMeDpVj27JFy37sn6wsoscIkjOWlvHihW/ohmCIiFc1Q5SIF
E53t0ajvqNsTXy/PXSYUYP2fZ2x979BVepiKfkQSVq6UjLT+nT2s/TPz8akO9P/P
rMUHHIR4MehyL34f+uZ9n+oQbyoEXO9L13lqAd99HqpKABxGMVptwaGRvzWzYQ+c
qc0JlTmvj2HeR7oYMrMeMbZpuFBhFPqeCQ21TyxBRg5byKmbe1T92OAcHZucSlAT
jYWPzn1/kePuvw6VlvesrZ5FczBOJcVLfEVZ9s0QgXOOFLKTb3f9FVrSswELzBg4
GnOiv5e5gUwQqG01QUnz4kGARiG3kCTxm7Yqigm3Te94tkgy2pKsUF49yn4puuqQ
vdiX6w2keeSbJK4OqHy8g0hPFh5lzfIS12MqDolkgtHvjY5rYhvljHlcyqeqeo5c
NeJcMA8SeUjalk2S8QrJ1p0Au8exq35TfuUa9tXEgWRgOQ/oXdBwhviuUg57RlJi
zEcizrRBftiRUHKREw+HOsoYo/K6rL9Phj+/2AFDqWbhKlSkyewlbCZV7/wlUI+C
xaNJg+I/j9NpLtStACbLsLg1MvwaKvgqRdUabw3I4HHLo1fdD0E5tAKBW+GDSaFx
8XG/TlYSWPs5uCiN0YaXbQHOiimgho7UeC8fVfp5HxM2yIRULpOW2PR6oLTGQeWb
8aQiy5GxFGkxWPb9N8Y+L6FIbQLCZonratFizF+MNL79nBpKdf/+jLG+tXoXBPtq
3FjFRbKPDc2uc6XfnmApkeTtcKP/4BzwP0L2mXwQqOEu05Mylf6WP5qy0eOoxLQh
0jxX0fmlIc9Ox6BYHYswFObXhHccYjVsGdC9vTzKT3lgKgv5FXEb4xYgY3D+9Eg+
GePcUCq0lAlpA8tbP61os2tDjTBXhENLzPt/DQzYz+5cnxfJT8zSwKvfkt1zFB3Q
ZcW+1JJKjmqZ1fuVRJeyNopVkuHOwp9R6RwapLr40SNwXRvXITPeMjbaH7XIbkMV
v9CPSRPynLS7cqysiHI9gy79oG6pZjK+8N8kWc2hMEW9Bq6fzr3YYu0jH+JblaWQ
z3cb9x3X1ygnWKrGA/EZcEK+ePyF+VDFoz6V6lGQfbn1YSEOdn94R+NOx/4GhG/8
l+AH+PRC5oUyZ94Lvy4Q1jRBVOaSYPmZnrbXjpnxlyy1R65OpG9PbfxL1M3Ztke3
q35JqLqZ6JgCLrbuCboRICimRByddlj+A1OPniMaeDQmHkz6XMR4FrUfb1a3Jg0s
EnpLmbBxGWOdcPC1rmVs/4HBqoLM5uRoNp5lKyoR+lx2WRLuq9jvgYL9q54A5oru
wnvEeiR6ogaV0qJkw1BdWsG91Dg8mrzOR5R6uJ7H0NEOAR8hHbPPAiT8acWQhzg5
TAXb4TJHcHbGDAfPh2ExtZhBRtff8VNbNqwB/0v4Ab53i5cor/1P0OcYcc/qKMmf
zZAZy7fev7sJSXdzNvR2hdE8g3vL0ao5VNzHPHxxKVIteY6H5pyyRVMwiSN5QXJ9
ywkzBt2ykWjuUVgfm6IeVd2Sx9eOcRsvk5S+21muNQf1RcIn0R4XPwYBrzUdjODg
WqWLXfbmqVC4KBE+ra47KiBjlg7VHGNO4nxvXFThcLZaiK2F1wH9bV97nV59GhBV
JTMGeJcD6P/08xwkM7S9Zdx0AYCLseLABb4ZtUd/nvYUISfFGRC+MAsPcwYTU3MQ
QPPB5CYrpMn0yrGWicELTQdHR9F90Y2MvRWFbgIIe7iMo4QJbVSMDyY1qkCBL101
K1pJmn+6uK2TxjoAzPHzWYjF+8cSSU3frsaOldcyZPV8e1GaHEYC4FOVqdfFp8ZG
fA9JizNS6UgHZ0HpVOL6uzqLqx4WHOTmQx3fDxLfEJBdLdZp68zmrTqsszJzQ0Gj
USKNVyN0lGRCpkSdmIkauSi4fuEmbUqJps4Qqm1h7rK2UH7DdShZAhgQVw+lRn5j
5zOw3npQ8eug3P/WXZ7wxYE2mo5jMY3gecftcGDCxZd/MiM22/QxV5ygrg4BgV4A
GR8AaGFZ5Zyrzhv85E1LlkVanzM4SgdqHT0/LxxNh5aEMD6NoHuyaUC+1g57IXTW
VCY6Zug/f923hgqTJ/NaWr0HLDqjvmPG0HbobtaAhC2tJ8OscQqN++nuJ2sMWUDk
Lj8alqTNWJQxZROdlBS1o6OQunc7dDw5HuR/2aqwvTf15KzmCCCAoCZuhcKO9Tw4
JP1bmh97zeVTdBB93/Ocm2gNQtjXgZebmFOxZTVD5pCf2KU0lifFZdlFQ8oGZsLo
wDU3jeBJUFdKXbzQrC2OAtICcRS2LlCKKybovsuuKmAzfrI4l3UWvBC54UBKHk0Y
NRmbRCBqqgofZXTU0dXnQJQPKMeRVsrx4zqmssnLf2zPuY4K5IzSGIR64mEJB097
12fJSKZdjqGu5gnSBHvPwjbM/XU41lfiL6JMMV6A7m2GJeIIwn9GccnR/zl/1yC4
N67JlF27h6pmXpsMHtrP08j1tKTfrEy3XmR7nV69f/1d+z8Ig00l17D2QT8BfPN4
mXZEK7Ow3iNnC23yDTrG28bWblwUULjrXWGW7v9cN9JBGIcKP+nSz6Iu8UK9SG6z
+w1N4vZk+S1YLVMYQ33tvxdCMOaa7egixKHiarTyGK1VpIHvnS+uJtRQwAdH9ZAm
tutdj9UrnDoaD+ZP3cOEM4+4v7BXauBILUgt+vNiy7vyhXWnZ/a9o/b3r0wE2YPp
cstPw/Yb+HMOliTgSPW/P0iITAMSNSEbrnlgNee88DFX+qdrk8wMoF0uO7pOmygi
61rFZ2WPmeMNl5xzAVbvtjJClR6d6gZfCnYzXDyDzwSVNjdmG+4ZL5D8t0WWB/qS
v8qcV+U1Vigu/Tfonol+PgoRxkmcgj6j9+O9D6au+ZVsBpnmFM/nc5q+Q4gmVBx4
8RlOxPfubrpuGZyb1Ytc99lkoiuMQIYdB7KLAu3jzKiDYGf8WwBRqCdvOzQYDhiM
bRQdATQbKe/MlOLEP4G89Eyo7hZgmARpZ6fVffDdg8a3QqmCdMWvnBy8YTxR/bb6
HArHSwCQ61OYhnBTqMB1PBRIbmCnC2fRtoeLsY54IC8XG6L1s3qY5VvRJgU+EK6Y
bcH9WohGstqB5+qjXJbEeoESaY3nOjFFPv1AKuf6pY+A2h7YH77BW8aFGUsGmUpG
RG5H8G49TRWkU7Nf8zYtcs9LM+ETLULQzF+V6CPPrGj71EOlQaxK6bwncCiftPWC
CeeXv/FsNANaUemhiWnZFFb+owkroZlBB9QRJLzRi0hPSkug+UGzLB/OkXKd3g88
sG6F5FVUVAagcEHG7NQL32lMyM6KF0hSM/DLhUMTCuspoVdNvIWEkoT1nUydK9NN
9ihYLj1k/oFFhvTXvSLxn1yNQ2RW11UUJwUNVNjcIMO1cyvn1sE5H1IpyYuqk2Rb
LZByj++VtlES3Ok5/ddv4TyBJ/oNRlLEkZDtMFT8vbrPcz9/URSKoVRgLhsM6X35
j8JgcDsuLPVCcJXfmem4WiQ5IU45f7v9Wcbbc8K30KUfv2EjqGtJMm0NaunHERhN
3Z/onHyZSSTbZUFXBqH3y8QBPhb07jg8CeOpdUvXXIa9x/UtTcGoHwn8chb4rhwr
Jh/5GC7EJC8LRsE38gRxCLrYdVYy+T9fbyCzywDy/t99OqcnaIj2c3zRvF9qWb94
i/m2RygGXvjJomHFbxQWYLEa7vJG9Ju8BrEqkEBKEBDiHASyqZuJAFBvTiM1N694
MCPRQWG0Rn8uuUCE5x65IHn66K8AGP4kjCyTlTtPZwfUrYivsXlKq4VL2yYY9+Rc
tUfjOjjAntYg7mth369lLxRjZXP7s2YfEhBkp4LZv7hTcAWgQeyA1IVZPuS6v8zA
fZ6duha7G5k5fGkJ8NNwEzLR0Nlo717Bwc80mpmFKwmOJG6iyDgMe9uADWxDZgJl
gLKtInoUkINwUBJkQaG36R0v+yVbaxkZiQ7TqPM8O+El0Krn8/j8HQfei1+vaE/q
8LBlAgs5T22i87MjIEQHlOFRWgb4WekEze8xOaeCqoZ5krr4137kBY4xce7YLmNz
lyp+SV3L24u7DxxRy8VFKXn7VKqzwk/Ewv825HEc3UhSX3KjhH2WqMEloX5/u41D
1ggePK2/uv4wacDK2WcMgtFjAfoIY/RVDUlyz1fTKqge7vEn79qhIWmdD49ZAP71
jkb8pELmBJ0+tYH3Mcv+v2hYiG6pepf5DNFpaXrRAlRA1C5mBJjb7wb8oRT6IwVG
IdhpPN3iLN3EL3L9oq0Jt2O4eSGBBvqzPxSCnZLlyYFiTXA11/7RdYADmbd0JBH+
BNs5IZdHBnHZK2XxTe5piDsSdjTb7nQb6h6QZcte+mEhoBJxWgFYkvckfs0dHhLo
mUDX9AtSYZnMKHSZyZVmxbQUbtIriB+XEP9Y/yL766v2/y6El5Nkps4m1ig71EZi
HymwQcvUXf1FU6RyzmtdFnDi3k5a9/1vQAfwgQZPPtSqhb/Dr7sZJ1tXbKOkUot+
RNas1hbI6Tg6XyYaZYYRg88LF/ka5aHY+5FF95KOZ8m9fY7YSO+XkVj3MkyeaJk2
pX+KEWrqwuzpaidm9tU5HxjXZTS6JK4UY79UT6OyrbAIyLn/muPSqIWEIX8FGzfW
xHE+/z8iQlws+CpCd/b4gpQdFyWrU7kNYEzCpWeG4OkZmkKg3pYUl6DRXWjIJa8s
akDsm+Hds33Z+y3T1HDZSTOXUvtpaNMBwz75ir6UG98PRFZVVSA298cX/AtBdtrP
xIoSgakcYlx3NiFA6YcTvXJkJfmeH+lXrC3+M/K+7rD9Q60RKMYQJ2eAyM7SG9eI
74INFyvvI7bmO2UgaBUmjntK1xrGtqwIyxoJsKP3wmw8ItdvOjy1ocdGWRV+rbb8
xATH2V2uk8NT4Iz9NzruxrdajkORyhuXsgtO3u8lBFBFW+suAXg4HcISoStDW3Mx
c7/hnWBHqcilBtb4py7c7EONSF8Wm+5ZlnW2AV8nSnYDYD1C+8wpUCxjLn/7yhKr
5G40SiTb/CHmwVer8thPZ6I8iuQcbLtRxAaGZKoIUtWdkOJy1hat3CzhQDT61Gky
OnwGbgHI5FGHbQ4WXGb7md1bvXhOlW7KIaL/bYzHltHiARE+iY6Gh9PmCrcG/cwT
LaQRTdzUGmrKRxTOTLxMiLHKaf/Vg7oV8S7k52beb4x88obzRABhqAAq6qDaDPJm
FPnFbcSGEOY2OE0R1E1+zmjMcUz9k3au8WKaTpWYKWCWBDMoOPQpWjhYSbryA4HW
7po0AV7RBap4dLhvLeFQ8aruAyi32lMxjgJPbwikbVJp8cW6Xv8hoNfj1JdWeBN2
R/QZKlOvVLZcVvzJlolilo141QZ9bFYSGrfIMi0K4fnYn5Gl1i/yXTg7nn3y39K+
qt3EaE0zecraZhrx7ettKsHCP6cPYz4AAxSCef9jGYRObr4YG6ZzOtlS1IS4k8Ms
eBw6oN6Ukb9vDgPRzGSY88ULNaIBxPshF3N/El+h13P/PpPL3c9dnmdu20z/8ybX
x7hecgQD2v5ZwqcxjesiCBGaUqMm2O1LKJBtePQYM/WA9F5suaQQUBuokV0MEXjC
36/hnHCW24QlMP1+8CDxjx0debcbpIR9TyTAEivKfmh+/qy9iif6A/vJkzXvREIg
7VbB/XeCxbP0XJFIc0C+xx9qn6pbN89flHrEbfZ+hVQ1c8KQuVVtvWNrH2N3jRDQ
EepTAlf1PSsG+wRnkRVPkoIDBwfoHfHv/YGYSl2K2rYwTorKXUBzTqLoWE/M+NrT
cTeVG6SkMUx1xnkmdc1ptwFPpj0nPSTb8M30JhjJsunBUG9Jrh5HE3s7h/nGvfXi
BX1fL7i7RUMMz2rqxLQCo80mrHrmyWVhbnbPaLUKraJ0LbKPHkO+Lia2A7PnhuJ9
719nTbcDpVetlvmEMIPBL6nKKDR/OeA9xGFp9IOu8GdF1j/KwfCsHdv/0lJEWXVg
BMa3yI/Ry5AmujUAnL1S5GbpwMnD72hTIX14Jd+w9ItiNxvH5XXPJRnquFZudTGx
alW68DKHIQvFv0UrsX/T1fV/2Yc56dipx86IMpx2CfPIwPGLCTDtQmBUYn/YLDlm
QXuBTp0oJRB335E6u3xu8HN2nkdISPhqEVqYD6/Kru4fwZPMGyUyIFUkNL2183e8
tnPOHDSrKZL9aGjBAozL57ZVNsBQ+QDx88Kq8lHdWZxskyKpAHp1DONmaCkzwU6H
BiLHiXGSf4/DSWfRF5wSsKR94St3HE0PMhhvgv8kPIkBbNcughNBYpn3aGunu1sA
0QFmCuSQOQC3r9NXSQVZR9Vr2Iw4HCoffrkyKfHYl0binO/U9WJXTADyLgxu/MC2
QFARHN4ac3G9FsQ5H/i9hStJSClZvyv7HUPR3HQuw6iIu+gF7tnaW4+4IulC9hob
M4RhQP02w/NumgXp9DESprJh/xqN0QiPqOZjjinpMdyLYKDWPNUnvEZdvzA3UwkT
FWK1q1Dh816JER1S6SdR8H64FcnjKdF0kklORCTz0ugqUJNnqQ1EqIu7rAhuin5X
Ewi3PTGvO8d02vkq2cXUXCDxaS66pUGIAN3EYZdWG3+qZXxz/dfHlE76BqfIruOf
TxAFxwiKbvBSonHCT+FZMvsyxj6M03hAVO+g51EsFkBCNvUh2OsjGNXxHnxO2HiD
l1G2/XhMh/UkjD6ArPc18SxAnlX/AzfpgSfRCY2qhyds1bvm300S6zgS3dARWBIS
SeArUHiE2iXZ/iHFsWD6YUscMcFJXX203FG8qE43GXmCWfojhpFMMEKED8p9eBJI
4v9Ek61aWJmAMu9GO2nbj/evdNKEGzqIX63A4J/hbRpueSiKB+7D7TPb57tslhbO
whIpQBsAqOfole3NAhchL9JpZqX6nSbMtBkFyyTbD6QOSz/3OKijoCD1dCuYEUBD
PlQ0iUGibm1NSY5gDyh99SIxxjLIOmMT1V5E9HWQer2lQMMY797vBo5Dzc7skvCc
RPp/c3liCK95EL3KiZFRWJi1x3wZYlMXNzqT3D98q5T5/AeUPSwu86SBWfALRjUs
l3ULVae2oSJmVLf5bbiG6pBhUZk05RcwMmbtZGVKDCVVVPh/zTI8iM3A7XM+Y1D3
VCwwRVXPVrXtoeuhmVAUjoFbLGMa7WOkGWrXTjJTii8V3YQDaX8VPPShmgvGh6u7
pklVuIyG7fiY9FmnJpGZCXZnXa0asgu/iF4VWVRXWDHPXRyKh0f01e+69uzaPMGU
uHH1E4dCuq30yHm82pCIZk1sIyPtZQng5wz7+++HocNDjxC9VncHtf1Hp18JO1yx
SFlZltgkD6qMMMjVoGddbgfuOcpnEjAD+ZUHHipWhV7DgWT8L6JjChoonlMHsq1n
3WjytKdMjwo5VcAiTGzfQWgage4oU2mERuBh8V+PkomTtHt06L/Lkva6rP0teHnK
UK/7PskoPTe/PDgL71gdFt3bkV2ch2tCofQFAfMIAVZEhyQx6Uzs6W/7tTtwW4+A
jCDyLsH0gLbFwerRJJ3UqRhCA3tvu9B3+kq1WnjmBf7JfV+YP1xu6TPgNnYKFDZb
eSlC3efz9Z0n81eP3QRPne8mdm5koemtY8nBHQitqJmGyogrdyaMsAZSlMvncemZ
I5StsxBM3XyzBADAyAXGkVGnSEKii/b0DsQoeKwCfqBCK7V+m8vLNqxUFZrCFKza
AnIng34b5T65QRtYra0SynJf8UrSGU0tErBnXnPa1mPTwXjkUemwlFlNwJzMohwc
OzLVE9Bg7v/5q4sR7xAoSOu3PYof8crswHYnc2v4DjfbTSHlPDsiBnCIhrtKgLG2
uAFn/eswex69V/YhgxOczZ9nOrgCV2zFJ1D7ajqhQhIZIJsA2W2sEvq/bZYnGhX1
5FJHkIFILkZjQ9t1p9rhl0Y+bzvtVysymoQ92Qx0xtY2EFEnZqKqjBy6YtTbAY9u
iTmfHnpvpC7JJk0+PoUxjs7lm9K9eAi6J4AW1klopeFgkIDpE4sZDA0zbb1AlGIR
AJ4d4+WkaHXLbuhwn3xurLfztXwbYnFzjDPfKB5+6BxxymwXi/vokJR2M1H5gFeo
wVkirCSgKe9MB9CmCPdZuP2LYnRB63dxpdi8OxwuVaeB45t3peL5jZHD906W9WLb
z5Zs7+UPQqqlEgG4UllwHxJSv1xhYTzQWt7U18iAgp9mdUPjKD2TaXpJB6q9OGqS
YjLs2ZZDAVgVM7Ulr1YF4hfBOxIN0Fu+hOv5QJUVUxNOjnCrW9YE4HCtmVUBKaWd
Q0WC+eK2X3P/ynkMCCw0j/woyXfmC4kwDim4lyfZelxfi2ZFvRmU0SZrlxFt3ssn
QsVR9Pz/W5N4TnXngG9lYX/d/Ifongf2JBx5iHaHjDiVJnP3KFqnFfZ3+m5PT2VA
RDDzvAVPC6x3lxQtXgkExjCOsVR+8+ddS0fIzDaRlOBj1pJEd9/zgk2LCxBR25Xw
Cf1dyHZe7UJMXr7/EP1XrWKyvCdG22NC8CrItnYZTmc8vzrkoDK3NVNujlKgX9Z/
gU93BBEpCBIp59YvUhnDPGpQyPqXtAjyT5o0Dd0ST+VzljixloBPa0k4RPFLkiEN
pEVSdNIoBqzWO0vrIqMQqw6DzHn6ykyERA1gltEqlNhtxfeg2Ehc04RbPXVxjDD0
2oWOYfgGf5Mg0ScH78cwR2j2K4ApW+pV4izk9qqqKSIWucFyyIKZzI9hFtawuzda
Uklj1SH4Lz81ggF9dKNcxkLpOs6jSJfDeGZQ4RJxOKiPoI3QoQMK6IXGby2SWmSX
XKf16BmjRL1SyiM9jtbtdr/t2K9ZEZ4ysq+C6OhIakgXULm6yGnmGKx2MAl2m573
0srDZcjxPlvRRkN7ZB5HKDpyzbGHLdwzNdY3Do54cdgsv/S/A3Mxv1EMVy9w0LkA
YVqKFj9h5uCrnsfJLD+9hKkqkoA3WaQQfmajCqXA0pGDjRoTaxiSCApEmykznPD7
tViKV4S7ZqWPD/UabhjgVBcoqMK7oenRiF9vCaMgFZGmP5BSWrX5zdV2+VRReXfe
CrX/Nwo3r1isqrQLPNBDV/d5++W6UsxGPspptkJ1b+mLe0w3U/6AT33sT+B8eqtD
Q9KWTS+yK4R7vuMGjHD3BckDC6T6oTBvxkUvUxUz/OgHbEkr/bEIhbDlI/5T4tkB
RRe19L57guqc8/GUDXEyyJri+CGe/W8s40SMlFtD1MGBmw3EkhKUGuImMzJtCPor
gz/EZoPdsbq6Q15dookKAXe5eOAR0m62oXyNXMJiSQC5vyPAnyK6GI7Nc38CBetn
MCvmUKSCOaFKyqiBYnzetyVmgLef/yS9FflGIhn9VuIApg72G+tSmrC9A23OLB9e
o6ZN3/yeXviUA/rqM+F33S5C+SxsCPa0pkcqv8oaJ7fPwizaf9nQ0Gmoc769vWlz
Jd31/YOS874V09EximiD+xy+ByEYiL+Q4RqcAaCdsaluxoY/6ZRmr82dpoUx2uMb
GRie002/Gkgx5nCZCW5Q9ENErzwc8H8x2i2rx/SsDRQOdEvSlk7Zcqlu8H2W4m5N
`pragma protect end_protected
