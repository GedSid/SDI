// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:38 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pHbHEfKEiewQUYpf53bMYWcBfxm24kMpWQZWFch0399Rq9xTHhjrKCCLbSZJZo7B
IqcxZIYsiB4nyx3hcBFOrjeBOv/ba0LTvJT2xrBFrS/+QjIEAc4u8t9Q99F46fH5
05Buh/HVHBIZFjsoRYDIjYBzlm6MAKOW5SU0KK+hydM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9840)
8hPxWQDzO8yAW/kHyQeCYCHtc6fUK6kNZcD6AyUsay8A9wSPHi6RpxLHjwnkjiZO
eq8jVV12hHsHoFXZ3Ev9GolmEnAx09JEizHtqWJSzpKfwxsA8u/NhezSM0Yeax56
S8oS6U6rnxEmnC2E1H55UKn9J7r49/KuDw/N8eyFsP/fAW2CWURXw+0P3lJ2bgzU
Bk5uUTEr4peLWz2SQAjTtI652qRoFSDYScNVpSUyINlzfMn9mNo24Ols/g9F1P4o
q2d5NbSpxSuly8CgD+BgvR4FCdpFCBHVTFkbiUFUifBDiqohkBOFwQETpb68Rl+T
cDXzE9EEDCG5U7ZD/qb7tPQn4/ABeX3HCfVgtLNRt6WNcUzlm8do+9aMqzXniIeb
YNIiIKXHWMJBZlX/uobHNtu01p+yIVvsYgpgzyqgWRYTcIIH12f5yxrkSD9DyyKp
T06i5q71vGdeMIms0Yz0os6mlkGTiudl9yFPZ/y2qzzzd67s/XaTWmYOgGCtbQ2F
CCvhII1cDm/AMHaRs5vxL7sGIRIw4TXeW1cgeSO/oOlYmciIx3r1itICgmRhzXek
xTzNI8KzkoFAGB9GBVlRod7V+DfYqhd3tExtaV3+hRw/XlmdAeXSFQd+n75Q7yoz
fECOp3pHopTjWHPzGWzqe/pZn3zSW+4Ji8Lvc2DLPrfLvYGx2TJhQzGOOuwMwQ6F
X9uUYOMedITrAjeqviLPu6sc5EfyWSBwkEHivWMiV1wqV0s8R7C0hw2kuMJZifH6
lh2zaa8ujoh9t3qBi50Sqs11XuTpcKZQHlNnHMxgdaVW3MFWWl7COWIgN+jx8ZYq
pqOjDUEjsOhbljPLu9DE3PD30GkG9mE8Ghq1GPePupwgEPeTRVs7fPA60IScL0Oh
q86kEGKYaNx9oQKypavGl2KK6wAQyua3NY01amVwLThBSpSlEf1XupUjC+EPiTdU
LoaWMX1uFMPcWAJgaYNcMzlwdpOg24vB8ecbCaPsDQlCWQ6q3hYEJfOiBf3bbfV+
+pfoMIQ7CCH1O1l2IFiEA0CpfruzQdXisYY10wYLNmt2AeDqPexS1wx0i+JCv26r
oFSA/mUbAqZl7uA12vZgRszWw76f6Ecv5pX6fZROCY5CFrnjdc1foLU8fB/8UqRP
NIgrGzxeI3mtkaGRW3Q6sV3dIqPJKpzYQTaGJvx1RMFsoJPbiqazPwiv5Hxy9SkA
0lnsOQBAV7NMoo26WikkIyXz5VlUBqt1kz3csdSV4EynHrM64TBP+04kY07HxTUg
2C1tZD+BsnuHSfrm5t/z2ckyOjfepLPLCuzPVNYlMM0fYPUSNvWUeWHADJNqIdHq
XhXM5Bgj9nynfdwfGxgsbonzSOot9etgNVXo/e+iid45PXGg+EMnCVLjpZbodc73
8HG8/sqYKPLQPamXELFJPOZ2MEHUS2XJDkbQbssK+gU5kdSV3YfDWdaOS8Mj2APE
z5CIP5HGdf99hM+tlXB06PipMUx9M7hqT2z6J27Cr0hC2cKjXNuRSgirnOEra9yz
qflA/WbU6/n2SuVl4XwHQtuAnR8Wx6e4LXr+kN7SIPPepE1zPoj4EWvm85iFZ511
7Deko7p98OVp9vER2FmsRPWaCPm1GHVOiOcj+j/yyPAHC7jh5nvLkpYWHQmzEoii
cxogcUCC5rKkw/H4SCNDYj3CfPAiT7DMMOuMBho85uxMZPGjO6DMNOtqr9HkgARF
wREcuo41LpbJdGTx9ZW5PHnbvLeiSnAGK3wdqVKx1Y/P1wHUJLqQNAFijDBT62rq
O8RvYahy+WRtgQ15+UPVuhX8T7gWbJbsg7HceNqiR+dE9aIXepYv/YqoO1MGf3qr
07cL/VRK5EcKk+zaV72wxPOyBw9oyWXP7plD3D93ZkzyV4aB+LoPmVL+3dRWmGoj
nzXtQSd2yuo2isX9MGwUFKjbZpQylYjySuHK8FqWX/FCeQQ3+VJWv3Bd2qa3UuhK
yJt9MjL4BNO0NsIUClmCLvTC1ngbFyxhtcZd9kxpk09N/ShK0TTAvrHg5tFib7Sg
P/8zSllOc+q0uvfUAd5bzlGTsQNyjFPzxT5x4iDl5xFtlFZorWdfzQD64E9Ywvbf
Ng4f25Apt4ZLXGnZVkGmncEK6/CvcUyE9JXXhwzqWDzWQv97Mkl6zydRWl7nq0aF
gCLUuRyW39O0CPibyzNk1DHFbogOYxSMHBlxbnE6GTRI2+Iw4+wfvTduOsZksbW0
zqi/ndGxILRBfsCSjgT2bzU+sLXMluz6nSG0yVj6b0sM2eFk8Vem0W1tQif7n4NR
6pOniWUVkzTt2uNwXg4/b+juVXlOwmH76F92vi9BIuqgukXSEpf9lHilodI4Zl43
TQl7UIs935MfatiSH7pFxxO65UUPz2I+7MQfZ4K2HZUnyiyK1ActvXaqZjyjo+ip
/lDlrf+jjIfIg6jJ9phozhUfmMW5gHhCtsISBm8rno7xEE37PuIPgBtHQhytnPZy
+K5WGQZO246NVbzZE0z/+QFGm9S7P8fJjE1v2w4tbNptkPhXZkEG1GDKfeRqOjms
xyceU/7X+L1a18Q/Nz+RT+l4Iqnlef9faT8MiEJ7WnaclpO/59lwLsZo2dbhgGkd
RPXx2b22y/eyaSAUzipyjnfqMbPPm00+H6B5ebxIwF0b65g/hawPeHOiJzNM8cd3
T+h3xc/Wn6ZjawtE9zpEiEsn92JvXTiIIs4GjK3kJNokrYRLOGQs340v/T9V4Amj
etXjbYboLScOjXYtX0HBsTkQr2zKz7CHWMW7ZhQnjmwvTph0IRQbD0YClfNr6xwq
HD1bxwnF3rz/9H0h3mz3tv7nWe24jmk+WnEX8QuLnBwUdqFOn6JWlxU2hDTKmkLm
3F/1zce62qjMd1YphJke0WYnCkYa6DUGJ7zdeI6eOyp0X8vvE1NnEmpu/qxdp5IL
CPhJYyUtkdJe5S77BV+y5fs5tz5w+ikX7BLEO/R9e+ZCFYYx0IRpAIHtJGlWny5J
jpY9bvS97Y0mwD7xiEWyghSUWfczeJpPfTd6msn/uQDP1qRXiTNtoua9RFBWnqiq
FuIz2Inm9ezK5QxM45ygLR/1HD6QL++dodFEcXaMHRVnqr7bwB21OdNi6x76kI7P
kw5BOsXoJ7HNOERYWUchwo9M2iuwuEXDfFRc1TlmJtuT1nyI+5VeA8Y46Dtvapir
1AM5VJFatALZN45NI9EtPkN6GN3lTD2uLmyo+viWo153N85bQMuD9eRq81voHAwU
iqG76ZRaxHwnt19FQbNTkbSbtYescf8StWNSf3RcPWVhQfgGqG65tCiAIjGUgCnc
dJ560/5vMitvgnmQJSAj8pvgkwusa8/p9bkzKkNSHZBspr0CrPcpH2MyW81cHiHN
t+EBn91HjoYB4OALutFw0Sqbu5+qfdPJpUnasRft9klppe6tTkHwVmx1FRdFWeOZ
6eLRvFERPXND2pYax59+UEIF+XfwkxgVW5DwDpbBPcO5ZB6iIBPXVYHLw2f7Vad7
4Is4LduJ+VPcR5fL8G2A3KcifdOP8M8TBpQbbB1cM/92wnfNmmAahwIaHZgQEgWC
VNiExHzGX9V30cZ1mdH9Udo7lku0HPF9VKy1hLRxERoTlx2e3BAilYLIylZbaqLJ
1eW4M3loE6QGRJNTTe/VCSu9i2hdAFNNaQpGZMKulF2D1IXf0TLMh2steqsaj6SD
4NN1crVwpGTgEVOxyhzmUWovcT4hl/FaSV2MlCTOLZ9SvxGhUTVK4LIMiY2bX1FA
WaC0uXYwfneQVT7aNm6s+vsXdXW9M226U/rPqFvaj7OO7Omc2xapYs/LJn/06qVd
KGaJv6lNbBL50IPt6f1pOI1onrFg9tx/i9pRTgX2D9IpRaVh3yxDJir1X+qsDESB
M0IeAAlzRURBCDS9So0lSyh64ZOiP7Fs0MP+x3OTGkevxTcWXYnKFAx4VQl7fkgr
K/8hVrC8S3EFBsnbJWQaWb1DXILYwKk6g5ZCIV4DhxHA8sjYLKM7GoN8AUNtmxFr
EdrPiB4av/F2cx6rBDVWVoq7mHsgwIksnIocd2hpBT3b4mw+g18hk/4a6UcoYLd+
L9btLmyrzdS+ep1Wk3dzuCwAV5VHq+bl6BN7SIVogLfaO8S5lXs8qmwEb0u+fcSv
YOPIUOJqmOiec6DztH3qRrVnW245pTjzn8MXSH78beGv7+uDKMFg2NTrXTAmTgkO
7amdLJ2Lt1BEg1xjLvpWqtSg5mvsQdkOmkVAQZ9RSfSfrkKRjXN57NuMHVq6oFm+
21wHmYwxGS04IQfo9ZnLzd1J2ZgkP/ineq4ePgqb3Hdcba0PajzRuxcKAj5apeJE
qAuvfWrPJYj1k7aczzRE56A3+EwzigBQMkjp/xroBCUfAk6zqpRLI5bl68kwMN08
UZd64gJ0mbUmwYd7a/u3VDBarQjfIUmEbqCtjeHvYshGSbwotgkeaU4U8VmFg613
DXxGLYRQbVtG6lOXFyDPnGqzXKSAuYLiaJecpZhGL/PEnLqr7/j3dnHp5pPifCCh
0cpZfAH57DAWysVIYUiYIGanbfyxzOfYrzGh+H5wJnenHnR/Z+WPHzJTLpCwGhej
aKaq1JpTo2XCO2aFnHK8s1Lxp+wOHfk/t+cQgjG+2ne06IPuN98xWfssXZiEJ7+w
L0RbuiBVpoSPBZoKUhIXpZOH7QcxrsSPNX2jNlcfFPoNnepdmDU7MxMzraJSIAZI
krTkM3pyfN5fjBcZJPipYOsw8VTEH5CnwZtQLNGZ3R7Z0qz8VzHA65of4YqMZf2B
KiBNfpY+z8qIzcjx5D80kcNM391b7VCROMXi1hFe3BQTUTy1GXaUtqWJzy3MJvV4
T1CBK5NxAJzuSI6Sx6z6M1VpCTzhtTVHCD94C88rUrxbzi+mTzxzwEUM1lD/U4Dg
yBnfqHWtWGefEhZiYG0r8kBfrDNm6l4bAogPn9LzniBpyoE14saN1oh6juPoqCqd
7Sbf2KBt0buGUhGxU0+Ty6a57Dixp4dUc2Z2QRwFd6771cfKOKGgxltnSq7zH5wS
vwHncLLFye8O0lnrhgLJx1cZ0QoFIKWqBxsRb4B7h4/tasQ4CNsWwchbR/dGv60p
atpb1FIk3qiZv1wOupVjkNRLb5xNLQGXm/FaZ82ylruJzrD1AcF2JatWgwkdSHns
cAwCw42jeOSSvuaUSOowKbNfbhR2CSOXID8/PDaf1Op+uOUW3Pb8xPISX3mOnG0d
6OpJtTDv483Cf4hPaftEbgoJWGGSydbCgLIL75yWmeuSywlT85nJP5Gdw/G75kiA
R3i1TP8OMyS3hEOEtWRYlKufyJVtMJX4u5+sLiEZXc1is17jWGg9tc9GtoMHaxzD
m3kGbNueWCxMZCTmT6Sd/f+reoiN2Rw3Bm+XRY235VPKz1D+sYgipkyeUGzoWeJL
aBRnZWqhpCNBwXnrXSF+Lg+4ghk7x4zgJfXtj3PPp3YgF9iS3V14qIReFvBfi9XT
B2VMasrbO9SIj+L508j06fNDRh/3qPTYoiXdeoK819Mt557MgFidFX02tGq2OINN
OGj8BXAUBb4DfIoEojlJa+3slOz0uHho81KoCzxp2QPeRJ0cdGeURzQTNLbFyXKb
pUEGGf0hH+P4d3RcODBn/F7drj1X/YtXlREGxxlET77B1mVe84W5gmuhJEz+1HHO
Knys7pE3BQ+hNjsl6Yn6fZRwrZO65sBx1KrRn2bNvZcOS7I64dN0oTrtS5dxTB/o
LaVPB5X+y2N5wd+fb1BTO5dz/V8fQDc7efa89P7uPUWFw6o8Gah2SfeHkjn8SGAe
ZpT6Y/Ibe4vSEhnwFBOoKgu9KPTFn1ttXYSLDSO+ye/WwU5HBKsUoWxhJfrRYqmv
s6xfgizTp2vGNw6sEQZnguvXGGQACO7KykSjbGXGNz304yyBUMnIckd1XN5GV19g
WtaIs7fCTKUqt+KbcRHDjQdJHhgw/jbZzoRLrw8UmAlk9NOvi2Dw/J3mMKxSaqpL
y5BxQAjxYYE/Gq43nJebaCQWL8vtWoG7gy5ehSc/HM/E70QLcJg2/0oPsuDX24O8
qiVZMrb1MtAIPBluf6RqHp/Sz10ajTAZcU/RJH29ooG7Qr4RxT+It/Ph/VqaSeed
HEA1k8TeeYAwMb4DEEp4w4K0qW9lUIzZhQh7NymbtxVsHftmSKW5DtI7+O5pRey4
SL9HlW81EO7OKvSMIwJR1UH8/f51nPXWZzzABBW0je3AuQ43a7VhmsaV8nwQBsBV
B7bGoWIt5tDobPn2xrYqva4/pl9RiNoXO4cy90/Uf+D5ivRAV5tNnP3yVTbXJ/oC
J2K+8kk/IPyaskmD4X8hDzhfCSYvK8CgDp4gK2mVYLW5rZZIfqcBA3cQB0yiIZB4
7mS8mcKHznLyp+O8J5nRxS5Z8ZKko6Zg5dZRZU6SwzSDfl4erO9LV5+aWQijX+Hr
H5+tJr4OpMLhxvM4NCa3CrkYACXUqGiY3oav4q/ScjKereAGgB5GNlPiGh7xl3Du
v8t1pXIPDhgRV6PBJhQc5BEK6Dfw7aiiSWwGyACkwg4B8yRVHiaq7YQ2+vFRGxx9
pA90+EbdPafSqs4SROK5h73nHcj/4ILtvePdx/YGP8Ts40z6M87QuAhxC1CmCXJg
A/unQRZNiHlvDtrzms4VDOFM41N/YqXSe8OY4jqMlZ7bAzT19lQFNLHEnvuOAD8b
0Da5d4+4GGXvfCbxItzAc6INCWSI1b8Xl3rda3NNwcDJ+G+Ce8HcNUDaKNtkn6jl
Y+VVhu33M8SXgcaDu4FuwphxvTw+UT5Vvt8+eg3IBAadQZBnelJUdeNoWG1+Hngl
LvPgrAPxmd39sfbEzJ3jZFqfg8obuH1K0pRVlova4qQELGW3ivowLoRzc3pOVAA1
brl/wMvWTKndF22n+cyyE6evLG28WtGBtDtcYNFUrG9/drYd2Mu3i7rE1Fb4O4wM
HVz5pc8uiXXt343mXlbpN3rq5mM5P9fvmqZMEOuDCSw7DUH1y0NcAAw+0h3GyoqS
FvDYp/td3dEOc2zyQqUwv66VzRhCKcfoAaiDsYkcaaHJeWUHDAkRGVzKXI2VD1Ks
xOGYX4O6ozwO8lJxlFRwNaW9orY4l2F6pVK09hEYx2dkLw7k5C+AuAp5oDiJGgAM
ojRqTmHalr6kn9j3JtUkynKPKPolklu16JXe5CoDthNCOGMNGvv38zxUBT8syxVN
1cpl9FlEGoDEerK4ravGKIMjLWXvf0ZV5L7AksX8GrD/cKICE3qeLZNzWcNVsYFV
ABiybB0MR2yIPv6bnpsp5a6w6bJid9IL1TO1IhxQhxpqSvJ4+Yioe9gMrKGsaRaw
+P/Nid1xp+cP6j57yMHcNRqwm5K6csbyaCzTIepVVsZpRehxI5iRR2bjx/2nhMCn
7R32Ns0FTmtNGeI4JxY0p9ZWNpnXRaZnP7LaXNbJHZ3PV6tvMS+orzUhp8stUoxZ
suyam3j/gtYfa10JP/HyD3+FPD3j3ujUd/IC0kqdoSKSeCG+jk6Dl9YV0yICogUg
pm/pR2fM7rC+Ttbz4E974z7HdSEZlDe4XZ6N2AeA7enbwUXaRle4yeJzO70/DyXi
nn6rQqgQWr05MgW6HEyLAYSHpeXyg0J5nQ8SZ4+KhPbFh8dqedui0R6XljN9WLOn
Y6/vzBi1nyLQfPet1vmQZD7HzAt9hx0g3rIbdFwPoofz20QDBMlnJFAWPj8GxgWR
Eb639VyEiRd1txsZfHCX64/QSnvi42OkNrIPHzFa831gj/DZ/K+C0iTDip26Qzac
QPNhx5htJOw4az1aTyQL2GjdboGmzgGdcdS83LNYgpKg0ex7n+liflhF6+k7wF0R
k1Z/HU7dz/pqv3M5ipcymxiM5j2FbR0Xj2VS3LRH6nuJgsGW/A+4atGMrpkVoZ30
YoSk6MZPWi+/16nEyevfeV3AL1VoP5Ot0BFjjgwUj6ydQhFxhSqkuvyFfbanzTF0
5KR1U3WLju5TJkdbnJtiSxvQRSz5qBgxeie58/0mKqsYBmcSFXZRMJfN4veoEj2p
TBp2zpxCrpZNERlYXSDAbbSPONbwKt8iuMeIBJt4nYftep/+OD+iMWnEHaz5dCDP
i2DFkqj1uYBnJYsD4RxNjcw6aaBhSNXCbnbafK6kZoKaluuZ1/T8Hwd34nEh7j8A
TTMQ5J8jUn3bJGwMmAQJ8NrVEtaY/42njJSvVRSDntkrfWsofHVYOg9E6WbcB2mT
py8LBxkLc2K6Bo+SLFH6joNIRWgfq1mbqtSEvKIV/fmIQWgM2HjRJpKk0N83E4gf
TE7/+bW0k4R7AwonfYa3JqtU+cg193O1oxBtt+mu5JeFsz1/i//1+v8m/jl5lBS6
0Es3lNzEvvnTz6qxLhtz/fW8sUBXaplAg5wLjBgkfT+jwZXSTYq8eGbFCabnIhJG
cNsZfD2nIVvKuhLMezd7f52fo2Tj1vTtsIwYZ9kzvdYWICmAbE4eS3v9O6DzF8aA
OBXIFdqQHRqVwgfcnXX6/jkaUKqNBSJxxQTLIYH0Ju713ZhzN6VuYDbNp5Ba0ZwU
HCaFF5/5vMklE6UCFbm/2Skl6Bhl4r84Tl/zTSfVvw+/bcxuyF34ntRqHdY6oUtD
RVkPGxvtsrHDONwzqqmr65oqbhiPx79kpqVyfTUFoH6mp9RGoFOUojd34x6g9Fwc
N4l3O0ibzPVqTRG03qsE8XarsVx6IdUnghR4t2KPRvp3a6YCnKjFIlkbMNqc9NG5
v4yASuv8s0kFCOYwmz60T8cHy31smM4y4E/c3pU0zuyG3Z0gLiiEd1Jxqsd55BJB
3i0UHZ6cAnVTjh0odLP6W8OtZ6hoF86qFeNyc0N96HhBM5YQCZHtjJLm+kQ/yZNu
3w64BrXkrh279n3n/OixP8eWwXXCJOUHC5RUkzgRiLasCk+Y8dKJSX8bGC11EWAL
H85ms3Y+6IMDhVJohwT2IsfSW/9RbL0WG0bRkFpixG9Y8TsyT+hLmSLPZxyte8HC
fFYZ/PRnOrHUwS9ew9QdD4SPxMRAgDxDvhXgtkFimPUiQTcjkRQFqd8vCCbNpU5G
LwabBLKfMqvoQ+R4bcSCOph4WvjtAc37dLBiDb8rGuLHdVcvfSVJhAD/MV0R6yqi
9M/YsBj2eyL54KOB8xGJCCZslIn9kzvV23dVOqxXeEzRzsAH8LF8/xeM4NWpKAsp
9D7mof9b80yMIw9GO+NWhgwPtSl94W0PbqJkg9YiajPEdvcbvlh5/zUJd8MYtCO+
Dy4AuuKekfkjWf9xITt8UtzUEI4JtKti3ugf7Y98RkRhnNniW1iR3ax9u2izuPsI
CHr1snB9eeIYO2w0XeydAVHnNNkK3oHdUFBBmKLtuV84YiSDUFjqQScnxeO8uulp
zlk5bFqF8rHNPlKxLWEZFX4IzpqNPIggtzvTm3q9VSRmYig7ulCXN4ESGRBhm7Cw
MmVOYRZ/n+ty27QGM6t0ng3WPALRlC9rbYOz0LhDB0o/JviAw2/E+unPQ8eKz06z
5yZhawX9kKZJEkAbOZjCWICL6yN1FdTAi1z+SP7CUfBEzqSTqFrQftvIOEyfJMGO
15vWMCTLJuQIP2k2+pCgHYRmSve/lvY62qK5dYEDO6HTNAqc7xNBmh0omZHqD120
1PbAGBdnLLymd2uQz4Fb7Xt0IS0wSSW65s+KQ/qgbAIRERj9T0lAFuQKxvHJDQXt
wfpRr2EOOwqNZSbC/HxFTtiqiVa3zfHEzcaHVYFWIXsGA8W+Yj51dC9pXAwofbTe
gZOMmXQ5TN7V6S7W65LFfVZt1CRITA9/WcD4OKxkmeGzOm0z+U/rzSXjL933Jz+3
YscQh8anpnzw5QwXfN4pgrhixpUqg8X5BKc8E1IX2LZ2KhZN+RSsufoiKDzaKbZw
uAOb3CPW6zPlZATPx8CPyYpZkK8rYVa8kp5rduFhRE9U0KLI8LLjg4yc6tirT90i
hbe3gvmPdprpsO5JlpDnE5HoJ/E0NTBlcEsiteWFarp6DILgjhvOmIrZ0Y6C6+QM
cKbQeB3GZKA1KKnVGYcPa095AWGW/r1gj85unX4C7iCJxGP8YFKzUIq5R/i11cRB
XA6kcsTHavjaaNB4z3YTLNnPgUQdLW31n75eM76GfmSEcylhjzjy/gRLvjFmEhXS
YXi0E6wRyVJeRgwd0S/AQZKdiybwKUaWF5OVTcNmX+Aotpf1wVlSK3mS46F2gjRy
hhzVeoJgPBmYkjxhtafkIxJgti6YtNgqny1cMDrl4WhWr8pS+ivTm3QnHnp2iU3J
BobNwkDezoKBuaF+pxw7sM4Z8aAUNpBCiW9yJwfd00lP7bpLzmP5uA1kvs2FrNZT
a61OEt1+yOm00lpbCLzp/M3utrMYAnQnduiERqgiY/JXzATITIrNrbLmb2hZC6TF
uKpvw9KF/cUfPq1cXAXMTZP0ItBzfWx1u3usJsIaTn/maW6QMFDlTtb8TLL+rt1N
PpFe0Ef6aKE9w1hPfv0bDdXP18SYu0wr0t8Xxo93eoqEY9i/MNilsD11z19hdWPI
lNjirklyNIVKIkVVbpdvZSm3E2ke5IwxYNxyPZu9W2wqzCgh92PU+0neVHb2Yzw4
sIRgEe7zkoNpg6XvYOzobdexXQH0nMmz1fnoh4bVVrzL/3rJasxmG6wlZCrJ95rY
v3OZwAHzKXkpWOskcdsgY/pNBvVCGK6Kxdz8s7NWY89N9Hiw2Ql+6YrYQeEFbJx+
WoUlKiPEovW85SoAQeH3LhnZpzhjp7hsL0vEenvDuwWIb6buXNly1eWwx4tIFsRT
m9JCinAxvXT0Ny7h7yhG3p7Oj7u4Vv1BKQlyLlYodbYhWjkA0HxP9DV3IUlkBsjg
nmaXplcZvX5zqrSECUn1W6nmkfB/aHWrPnxY/O4fUQx89b49vfzqoWzyidq+qBSZ
aelm0uBv8MWK9zdKQB+iR3ymnjQOP3g0qlwy82guVB0/YaZEzUshSeWE3WU3dmvq
Qpty+dpcErgkkFnypPbsMXiK3It1LziOVPdxiWdAOnrK588kw5MQKlHyVeoNO9uo
pkd2C71PHbML9hUbcBFcTfRBLvlinj+S+OA5Nnafm6LgPezYs5CyHtru6pMEA1yN
1Om2WLaj9hRWRSD091aPSL35jVjT6mbBHoB+gSljGYp1f6isyNERhFTRlH0ok/0z
Uj2u+eP/ZNtfETbXPhklxFi6/gQ9zIameUUk47+h9zobr0vRy0Rj7sPWg/JXTCqT
Fuj7tPjYbJUt+jAuOncWDqE1eGEx5n15bohfGb5qLSzCNj898aHOizKgzf8ShB66
QtHL3iTWflqJtek8e/DpGEBeSqE27Yevny6NCVMs+prs9ycSKbBGuyYLLAk/sotC
7qi1DS0F0apg9ziXXom8cCPoQs6VtT14om1dqXqM7+PuFUFSYaokUVf9Zy8ZM0g1
V9+jGfLq3HttKIXDU785PEaK/j3nM5IuEBsRPTMDVqUd5fCVu9VHNCc51hFD0gPz
G98kjcxOplwwm4RJT/Jv+5axGPGvEhd1uKpcvFdvXXYVTJzZudu5RdP7EWLdWY+c
wFnJHGnWSp50/eUPmDajR7FA6l6wpYAVtOUvKTMpYZ0PQi+a9Abd1U7/XobVmqRT
HCdx28aJG80P9E+w7QBblThsDzVgGcVtZO58nSXU4GhhM+gKGOS00IoDh+hsP3m6
l6uIVP3ngRebaHG1WY8aZ2T+kZGDj1KaUlXw/tP6jxfLkc+ZySf7go3xib0jPeJW
gOGNGPbHLGkh3uDNOJPSxd17cPSBgE7H3Ctt0194qZM9wRp0uNvs6ijQXGA3aW2G
g9MTCZ4ODE8CVl32jbyPaASBCoCaY60F9YQlcpi3lrVGfCpNj89jL46W+nUmcXwC
nwGKpq/VWbT/Nqx+FWaHT5Ii3gKp5/9g4Jwk9tyD55s6J89CvRJFMC3V35oZY/a3
DWFRdhvPkZHjHY3KX5u0PbUwXfjHxsZpVx0huq5lo9DkFVPAWs/OLguejcah+Nj/
30csJN4HPq7nm/h7n5FftE0kvfXncbikdVJyOILj/Y2Z3wbz+NQ3htAzmPSpcnu/
7wN3zJvQxj4nobO9PcPMdvmrfHryZdpc1uQrSRAxghXa5QBdgmyvlLJgjygyUrJ1
F1r3EvkL2LGVHfVc1Wf9/nJdNshZImAY7gkJIlxGMV9JDmK6lWLzrVIkf96vEBYz
QCtkF1PrR2TJCTeuVABOqip2tKKegsoo7UoFPxcRsqO1oG++ezreVa+cjyLMzT+0
//p7Z44vQt9dNGCIYGXcJPA6WHzeSbjtV00HgYKvk4S2wlNBRtZmsmFFRO400ltI
nhfyFyPjaI/g/DjrVVQ1aWRi8Bi+swuU/s+goztdNGIaBdg2pLgN6Jw4scE2WNL0
fw6CDOLreF2BwD992rTodxaOIMsCEMLnTdn9DvE/M2FNTUPDLDCRTNrwlOJ5ZjMO
+xZ5Geqkm9Wr8irpEFcyznb6BAjyHX5cH8D1jBI3oDqU0JyoOVmXJCYUzDIyrRT9
nVjId72UZcKjFwaiX8RXyBx3KI+axCY+5cNXXZdBkYecaHW9g/F+3dgF/TYatNHV
GhLKpCR1kdXusoeexgmceicy4qFbBcaotavt0KXEVTJx0oVdGVKPA80Prp1zz2El
ntfs64Ov0CCYk/XwOtxq1PzfhZAbWIF2tge6eLfUVOEx8NQOVPk8XWB479uRMNv5
cOQRUaQk+GIchqmFLOTSJDHzEtMw5HlzSmZ2nbum0lLADohEXC2Id2z14LILRt7+
27rJ2+v7UIb2aduuPCHFtkkF+5E+262sRZIiKuqLyiU7YZCdwLizkBTdD2PrxA55
m2JqRqaSIxInLFRzxi0vxyxuzt/LHYkFZU+Cr4HV4ncTHU9xGbUUaEwkl9ZC9lk/
EVqNhDxCunw6goxVVnKAHzexddLWeGD5Nd0j7QxsnO08HKuws4SHVBmyhsBAwheK
1eHRoEp2bKobI6EXa8ba8pSI5LOZ6DMr3rcs7+321DgMlu9dds1fzDX+rjxiDRPP
CM+y03PmrNaJ0CfldSGPRrXOybsyil/RdXXHDlKXKww5NDXGLt3/MmX/EUhxqIgm
`pragma protect end_protected
