// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:38 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
USQCVGUijnTyv5izgduaopime0VNNbRR3lDsDB0rL7eZ/AuJxFvXUaXkUuOsn3EA
PsMdkXg3GuwJnRpEw55m0qTP5mGx02aiG7Cx/Fje1cthEf++9+dGfK2j3P/YzC9d
hVNdmTP28y0L0tdfKDPSrxxMwVXrl6XMSUFtKiHve4Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11648)
qODWzN4TW0JcUrr4qpwGMgRp9MtZzFO0YmG7IH4XUTIk8KPTFOUzInecPzOy4gjK
cYVFmHW4mv+GiKwX/KwvcvtFRcoKZGsXdGUcWsFdBGacTzhztXk7Pn4rcKYwoqsG
R5Y9aCrCi/Yxvi+06VdjGF58xUCTnwwZWmY8VIoRSzX5GSBPH22ERu++jKG3+vyV
MzOlW+Ljk94l1D1NyD6fpjYbiAbVAo2XOzvtowjpPDW0OLXfqITJ5FTYBaB7wYB+
/0DoMhxSQYflojBXcRzKFU+AuZwpGClE5/Od0nJ1441cP5UWQlOZsJXMQyppneb1
APR4dWyVNCDIRIqBYnOnOm3XubbzPG3Frvnj5Bh8mfZD8+VIpWfYcpCjiBdcfYKY
lrV6b6JxQzBgAmYv64KWoXFTsrNd/KkNMqxJUQBOZdyPmvjsuPbccyy/fWAldc2D
xsz40oKZnadOBa25YgcrRV9Yyw32Vp8U9VzxBSVKD1M0ZPo9aLj/hH0STHgX/bFi
E3MyUjcYp1RL2Jm1VJ3QmyLrabUTLc7CqdEqIcPaSB+evLiwYtne2sQ2giCffM/5
JjVkTrhjTLTvsHQ9VSqC1maa5MvLN59YU099bQ6VSWfXv98zaR87pp/iYCuqJKMp
P9BqyPwfximpEXHl9MgfM1EmfA56e6NimtwVsJK5dORvFbDehDVkstNenQFmhkjk
hffr9iRRS4vxZJv2YGiEGAomzg0m5m/krmjF5L7SA9+zCiWPxZWoafxGEfa8iUc1
yq0CViZyLu68nIYZ3Ge2LKq0ISH8Uc6zgdde0np1YTxAbVxhcM279YQyTylBMx+/
xcvRe1QJA+xSVSNA3EOJLjF2cuUi21Z+mAbFFZVGu3j9o7mjcKgyEvlx8pwiqgUs
FpkVA8kWukB58ao2aKBdi5mxx12eRPzF4y3o0vga+cZtda4ecvr7/Cv5tE11TanJ
CTyXh+Zd/Q/60px27+O/xTjS+wu8V2c8kPp78jp2VNwE1o31Rm0jalIDp/LaoydL
QMcXCNDK0qVX3JssHx7Z9ZNjqBqje6yRgzM9+U76VBusFaj1q2Jerx5F4Ha65Up2
HlMVeo6GyIq/J8BMbUVvLJCxQsISVy8ZGbDipY5JUUOQTos65sQ2n+RsJ5s8OpJ/
Iqm2Rdj3g7i15Mrw38HXpt1haiKSOW2NIGTZp/+vLIF5JUwthzWJoY8f0WxlZsa5
NFT1eE/wjigOO/YBs7kcqjK8A5rSFHj4JPVr9XnWNsEsn6oBluG4scLmKHyjuZMK
YtJbDi35dFGdd5XWVk1mF7pPteKL5UQocWQIUBtkIIU7O+papca8TM0TvOXLoBDG
Nr1chnFaMybgxQpFbV+mFmv4LaCI7xKXZgS5ZevbwplR3muaoXCA4vkW7pwkrNy7
j/Q225PX+Xu/xHXEc6TFHO6k61fICBg3Um3hjTIBzgFwTeCRkLXIcHv0CKBz016s
Tz8P5EwPFbsxhR0W5GxFrmGpjK4+g2K/851ZrDFzNLy9mOPZTNT5C6MqkXeH0qcd
GxzgNDN65ELQOI1eBNTus32BOlxOfL2Up4+XgpZz/zY9qvTXBp82StJKs4Y94NI0
sDXJfrfys8uUIAVziLJIMm4sebkmngcLQFWKxk4u/GjFfcr49JECTvidLr1OCULg
DBfkKGIHeOcTezvTDqjkfqG6EGY1cG+lvu3Cw+ECMXMAsM8O0Obyqwh2zX+1JGom
t1axxzGeQjBgdU7BD+1K8CYhvAKtBWL+mLvbmWKKWSc+A+yewkncptfmUsCsk2Bd
Qy22nTobkJIoecwiiEkLiHJR4F8I6IVVpqJ3EESzlSS+QhBxoAwHFdwQTDUfkmm2
sOj02/fD2n5AmfJUUbo9ue6xXepgTrN31/+nweEMfqw9QqW/3IDRij/5V//NFIvB
OX5hW1r4V2WSm1934NrQGNzqyCBSHen427lXHn/qnAimb+CczS6ceHuXP/vfcavo
ST4v5nx+r7wS2UufdUYEp7+NBTDgmFPRx8Qv+J4VhHg057DOAsi9N0m9t6MotbyA
7ZxiEEdaNRNqjYH4BeVM+ORTr15NzvoV0PBnvl/fpbsg3mbODGVbhVinR0TF9Nfj
C7cXaYuRP0QT42fT/R4GZ+Wm0IKR0t+nbfCFjlLx1y6O2JsOM9WBLwP2Lx9a7AlM
93wi4cMfjZS4cAJUve8IfVWuYlzrhxY2VSBoJ1wMtByJ5YG3cv1dtLfkKgysOgtv
GqMmHlgGezuV/yiBkXzIKbalMOO6NEFT4KHljkPqdkLKrV4RZBVyQ4TlicxxpvNK
6M6/RU18HxbuSWwzm1Pj3RWvlWipwTfrr4OBpSen0xPfRE45J05boyrIg3BoxqnE
EApRvjAtCYQ27qSqWVX4SGPjzMj8WV9zNT5kTBSblyKsJjzjvCMBGZrEZ54euX7g
4qIFRQCVI9aq7Ho+2Zuiy5wjAHp8F41+ono7xrt1qzRBJAIvsMRZ0qxLTAFJy0Us
uXaJyYiBo+bdV07HFv0BU3skUOJ43wVQPRJ2LUAShdWiLXxwsjI+WT5913vwlmFK
T4rU03RDOoNJ5YorlDjIXaSTER35h5uM6KCCakog/n0ngms1A7BucywRFtEPZflk
4dIZyp5FLCKPvrSz4gPBkEEgN8/1VIKSsd+S970lzo4mRqs4fEmzCviYPTFCne2s
t6+VVVtVSPRd68klp48iQ+MmCXaTnpAwlNUIHMru306CqsHVZb7z7WGWL+Nefql5
ayhqgG6ssPSnsdD7FzFJnyqM7q1mqYiQV4Ht/NBXqQiU6KaVnaj3dOSudqsndE3d
tbsLpmfPzgHgJKXYwlMYioqo1U5fd5bLdyeCgiHBJz4KY6UURvTa8gmZD7GCqIl+
rigiWcYoytBDWc1POCuAwGbV+duwI2qOf6auH/uKdQkux10JzgBJfSeYc7ylLnRe
SRJWzdEkD4l3Hh+sM37y4k1x38jYzs/Zinexydm6OOpThbEPtlUfaAQ1VT1prcTc
28mhQBJe4Ys1uxVEnoJL2AmOp2a+YMHtCCatHzqpcMauw0yxYHfGGbPA7Xb9iY1Z
Bu5tXp5ZmMRr16EqYcXiMNRn063z5eRMyn8m33n9BvcIPOTudrwuqHIZz4eL99RK
rqPJrpGRNrto1iK4NhUYS93qk4718bzKryIgEmh1fOKEnRiixVXL/mUKFxA4Bo+q
f3tPmWRy1nqMPlWBnIUhLMaacooJ3e6XQwaAxu/NuJNoDrT1q2q9edtbi/VTvdJ6
JELhsWK7AvICGjxzK0KjOGhbCXydFDgv6UQ7xuTXCI9X2IyGXy3MtPTUTYnkWgl0
uWyIsLv5Ml3sWIs/mQliG9XSvf8s1e4ce89lowQIRtzeQeLjWaSQRdN3lpD4sWeG
2GRC4Rx1Rj4RVpRxBJu/eql+F+nTd0bUfp9ERGpAr/ym9goSG4nCgI21ntsJxQTN
YY2mawwKIObggOTIkwdVb0FLp2XySiL2c7qAm4Y0hxcDaPAy2qJDsNqWlAOok85a
pPXuVeKJKdgeb7qeq0XkAIBL6gAhs02glSnYt7rZvi58za6leTQYJ5BPyMq72oxs
LHvHuz6ylev/v6tVzGsOUlnT11dSYhkFlQg3SPCPs+n68V/YdPx/W5meG3wWzqQT
KC8flddrUWjD/nq7k/n6cfHaJCMH9I7HK162r29xUpeJ1y0snLYvRo9H9M6z8tVI
77NrLskFxo+8TInTapWJGTOzgUdPLRjtFF6SETaQ8+i/ToRVG/Bx17QwQ76vXEkT
38xKB1+Bc56DGHQGw4JUxEvB6j4i8Qv257mB7OURZynnaPifCtOWxOnFIELcZWF5
zXjU9tgBiezQRsO4TAmkUol7Bb5zKY89Gb1GwuxgkaMwnighhvq7CY5BbtHqk7Ep
38+gDjVANCL+JzOkViFBRrTk/CNeLLVc7105IdrJ/LerVsF7wfsGMM9xA/Aez/r7
6foY1e39GRUI8qDVFppxtQV8vwpvKDqa27x8I4JD8ZRyt8y9PeeumZgoA+AZDSVm
xCjvnTC8I7RxeMgJse8ms7b7xLDlXOxDrvH/n2ADSGioFBG14r3sblBYBDTnTQsD
OfXchhdFSV6WnrHKi2pvHE3JD1IYKi5s3APctVHPOSN7Pr8gG+B1eJbWb7n1U5yf
17lxpm2J6b6qDorM0okFQI/oc+Dzp23Ejc5rQSr9PjgHsRwTtP31IY5VZKGRC2iO
YLK6mC2L8tKWMLMUZlbQ5UIJSbm73hyWgmSdNJhc3pOcYp/TnowXq4MBDg1rTEvN
sSFdWoZQCNsNqdehxPi0e1CoUHUzyU4RgF1gMU3/T0NZtRoAt4EAmalPOrQYSt9Z
eg0lgfYuWnvsnsO7ToMl2TLbEuWV7qrKej6/J00S2dO4iRjkn/vtV7p57Y1E1kQp
gDtHfeCXHPDUj0yAFFK2COHCmF0ohc1MK6RqtaKWDMc4LhccUpS4fcScqHXuG5Rb
sWkaI8HEfFKx6uy7L4Oj4pI7m8IgD5i/48DSURUkqA7PEe1n9q+Ir3F7nW4B5GLO
Ef0Rf4AL227kgiHWdftiRnFSqLzpQPpdTiqZ/Sab4ZVw0v1XnEE7joKVSI36bNFc
w2qEr7Q+11oZyksmwzetWq/4KGMaOBbMDINr8VZG/C6ial0tLZ+QQZXVwh/G+EUk
lVz7UYSNR8HSuKjHqDstoJJezg0u41MaXL/P67asRf4u6J18sopIl2EY4HAX93eu
O1Bd/IddqmFvzrAdw6jEkSHq00BsgRRt+hREboeeLmLLZ9E/oKdsZCUja9FEL1No
dYpaVnEtwE33FHvUbis8+JtNH57pz4b+ay45JghsAmrVQOmzaOm8F4K94nllTChm
INYwbA4ixEQx83QEIkaLQr8EbmaOz6QTl6ImXKuGuZgzl5K2OOz+sietAggVB/oR
Yl+V5EmlFoVIwt9ftzofC3DwR0GBHwHiBJFpx1y+kctnc25eunJOOdimVx0llVm3
EwKFdfeCPYTDTfVaS2IbSHk7P0Qr966R8sV4l2lH3fBP+XekRzoOFyph4J0JVr7o
vtgh37Pr9vmTE0kZZaaJ5F0s4NIhQaTD+Pk5Y04DpnfzuoPOIRfMT5E0BjD9VPqp
pYcTW/CuAULtJv3HLypOfpf9p8AyjO7+e405C4yB9KRmsJZKgikNZ4GojPhWg/RA
pRLroFWyo/jJ87LGyQXCo9Dle3uFtGGtJfHTo7p3p/eWoP9MPO17iDTvU4GP1L2P
Yx+fJdzxX0gBvERSuXIGWoH38mQ0/8cB/aQquJqD++2fQ9AHy7sysvgMqWsTv1q/
K9wprjNqsXyxCWXeUJWtDymRQNKw3XFSkta6FFffRl5asJAjCvxh6qQOp4VqfCI3
29cNYs6NkXNhV+WudCRUf7N8CJZnr2ZFsBCUcoE5xLGDBAj8HebS1c3o6sNHpzPC
x3sT8ngZQLuPGxhq7g16MNm6Ml2DTYL9tdEr1NaajZuzf/pVWCH5J4bKdJWZc46m
RHpLjoXmF2P3u50SamBz04HxAgyIjrzzD7AnAbYtgingtMRAQ9z4YumTFMHxaF0n
3ku08DAAblA6/sPfSLpB5298B0S5lXoeVr0i1tyMwJ8hl3amSU+45b9NvfGlrwmI
lRW13jgof6BCNraQjiB0qWZEFjZhfUmSFUUaFL39NcRj98yx01EErk6YmR8spqeq
nhz9KPGyEVwNTfP9Pw/uCRaHzTS1mRHes/WweS/GxDfiryKL1baNg7KmGV5FebX+
AFJRL8ugSmLG5g5k/puE/jttcG9jOiFWWYJSyjy6FYggJyyw0kHI5zbx/Vt2T00D
0dnkxcMRU7RwdIB98fuwKYwxf8GqQncpn6o2MkYr57mw13wA9TDDuoAxVkkfq10L
2CwqIfpueIKLmsi3gOp7ahxhErxG8AhT5T1aliUarXqiGS00VaMsqytw5F/JBG/q
E3Q9CNTU36Xi/FMuqUCBfoMsjsTRSRJFxzZJpxy+oSTp69Bm88/6nHpbYFpXn3Pd
Igyo/akPbG1+U6Vuq9JUToKu4FAXmtfKs9MsvI45gzxRSBpMc1J0hh8RAznalD2D
g1ghvMdk2b9k+EsIt9jkjjcjid2dj1edsTHbsaierkRXxM7zj09U18U1IvBCDvD/
CGJ6u3sEhIQPESN21aP/mc2H9mg5H5MjXi0W6BMRngGVfzenCUX3e9Gj22HzDdvY
5O2vTBqEuNKVwD/RbhHz9S2oB4lUmcEvnwpTtueGiPn/ttqwO7jXmrJjE4Omfprj
1RJ4N/kprBo/WYXtoPxSdVEmF6+zTppCO+lOqNcJj+w8+5isQTac6MiqBnLmZZL+
se8Mp9YAdy9hYLIDG75oiBfBQIMcj4pEs36bxZCYeAkq9bylM9x9RwM/EuI2Vq53
AnABbUX7PoaKyhIy9dEiaHKR8jona8QiK7+KK5yXdwL09LRJVrmQ0eavovouN+6i
O6gzEnoxP7S/hGRFUF1r7gLXBkz3r77HSdZwEcgOBV9IWpuYxvLCctgZ277Qk1q0
zsU5E9uzTKX0d+tbUKkCcGukuK1XNpr9A7smsjZ+VKamm6Ua2O8CADExslosp9bX
jVssHKo/iJWpZf7nyvcCnRJZNGsTcquiwASZl8zIfPmioCErpFNqe96A1l0N38Ud
7vPfj9c5uxmG9Skh/bwBzTUNl9844UHCCEAx+1sXYHZFE1+pUw/c1hC2vacY1O2C
9j4fEu4JPsu50qewhhQydQOFOkYrPUCc36OU+jHoNnVjseccZGn94KwZZRciucUT
mmnAkaIKxggnkuTNEKWskj+HFUIca/qQSm6fnGdoYw3fFJZvYiwFjfJml7VhRrxE
Kg8g0rZjnJ3P7sHFyyDco5zEZ8VQncko1cNfPzvT5agdMMkokmlrAWcmL4/o7Idk
rXy1q3OALCYjgIdOIeCtU+8eiuGHqvH+vX9R8EVj2sRqMyRrpmA2s1fiK4gaUZcI
9PieGorqDdEcEYFSCHbMWyWHasKr9JYIwD+ciYRO7PTpq6kJfuDTOz3yGi2XLj/e
izWfupi+9ia0FT6+z/BZaKYwAm7XGR6uSKQQTTXvTWtT+0v7BWjQMDg0MJNpF9ls
+Xp/CWkQ3RdQBIpSFld2pdeUtVUqMvKzPVB3wxAhpEM/BU28bTd3p8WypPo/CKLW
T7D5PtPYpoxmU9+rmwDqC+BurhDA4nLwwHA8xdovwkZoDDwNi04xWuTny/devNNZ
HNu8h605DQbL4sXbdG35rvrB9vrKpWQMETXjh2vAQrI63mhzqptqgSTy7b1G1z5z
jG9RmC6e0gUnInv4VuYmEJwujn/hfD7NXjMRDTZC6DbowxnAGbISpy7tdE9/XjKb
TjWDzBNmPZRVp3g9AKvIYgizcOBDQLIpYbk6cpNTKasAkFGtsbcwL4d0qMB4nQcm
dTrGKz/ElW4ArTEQnFdj+C57TTxHFWu9z41uNhDIzSBxctW8caNZSp0BXOga4FOW
JhnIYGKnDoVSjJO/B4dizNBL/coQBlTDU+HfeKmUT6QVYuSFyw0UzQ46/eagC9x9
xTl5+anUxux3weNlwqu5SR04f1gqw3kkSGScGvCTtjKVGLDEu4ZAXXN+Sq2/TfeM
uBvdow/ryTgONTu1RG4/nupn6bKM9BNAe8ItSKabRKagKxFo0fADh+yUvqHyfhm2
R7iP18QuqBTddGZWOJDzxJ24LjAg+OM6Kyupa/Y2tGLXPmnmPjyj3nGZGz0qc3Fk
m62f2dF5Yi2b1WftvtSre7x0rHBGhR5BCcwRG5OJQpRGX1KIhSkMPuxVc2vsLhue
Y1Poc3GLIk6dYZ5l1u02jSFiZlE6e2PrTNg/DaHLqh3rI/zFwkrMQslz1/fYalZ4
kHAthDZAv8/pdiXA5PttBGz3ve23zchMAWtThcLDElJMYwTqbfpyCfuP2Lq91ctT
TqfKR2c3kuf6R86Xvz25tDw76oC9wGGSp1Yn9wzQCXzrOytolDWKJJycCo9/rmie
RDwoGsipxyftwWH3FhGoxaMxBlHuaSUKljk7n0Cfd0w9QR6xVDxgjzE2EA8RUumB
lNXmEgdRsqyhA8xxr1OrnoOHro/4Lat2uOdBYqYS5m0QTE1ndFLLbGzODRr+cudb
eCfCZb68Lzj2+VqQe9z3oMonAlbRsLvvB3ZgSqcJa5q4wKfz20CbB9+j5AHRcyD8
KTZMB/Q+mygXpjwVHtSEIC6AjscifGdXZW2UhOXPO1BfbN2M9e37zl08LUvxOh2H
Rd43jrUOPWJE4K/QqyiV3yvzWTernCVAKA8DbvtYNbMGwtPOaG1EbhMEtKBs8oQK
jQhj3tc6lHVVLOaWEoW5cPPXGE2eoNqI4Kyv80uj3pYIdR0Dpr5m2kXNnTzytE6c
TvOHJqYUyrAXB7wyjiM97dTCgFm/Mw5vGzWKCXSzZyfgsRKztr8vadEjm93mnyvT
1UKLKgZBEwHCtJVrBLI/iAsX+qzu6PYudi/f9hTc1R+eryZerS/m2xv2efPsyQ9J
fiUIsMfM0LUPdCMV7NjO7A70jS3xhxe2r7iWeCWmcKRfrIdg0g6hQ1szNBn0wZSm
7Xa8EmCXaqNAH57N6y4lAx+rx0Iy0xITuvZwXXiHavs6E/XlMis3TYU44usEOtbE
mCoGZWvgyK9gqwnrI/cAXqWk/wS+IRd2/gv7jXtM3fSyTp+ICfH4+Xr1oB6nPK5z
qPDYsV4/HbD7vQ7lTQT34vV+3zPxNooQGzLJtUIYJlQ51H6yJBItuJudB/RN8k2G
7u58gPA3bpcGSWpUJZIuqzIz3FpnJX8pwhWHRhup47KwOzv8VMJ39UEAIfqTmEuz
1bnvLYZTnpKuU87R+k3+vejc4rAb02zDU4ePlvpA4tx9kWG7cTGwlvVU0gW08zNY
cxkuJRe+BLk05FTz9yODWAr2hdOJ1MlRgjjhdcdqTi6KjS1dE7jib/WISiSEh2yo
Lo6UOPDrVtRvsFf40ROuNYY59ENbRB4wGZsH089uML9iVMW7qEo014RCVe8jFbln
HfyGrErCdQJfLnLNPuSvlHCi0YV2Rr+tR5D6X0VRlnzPFvT0tFlDFxG4EvzDIoaP
Ydouz6w3uz1B96Qq0x2fl6SIZyLaXtZj73NRfun4AUAoZU1mYZTWm6V+rm5xr6wF
eP3WN3jlpKMbxWNIBhkD78PGN5Tr2qn3FZI7UEW5jOaBRsHCcD9Fs7K616Gk88ie
3EQ/0s0cS1zSOmuibISA0kQRwhF3GNdj5pJW8PVvCSGHaBJjSxY84m8lM2EwCVtu
nKofB1uRcr9JBvyl18QjceAbNKj8NgBxT9yoVR1dtIybF/emOSiV2mNIubYMVneY
fp//8E7XD6Hpnp8KPAylqjoAA23A4VEO/LIQpfWJv5vRqMfAZRVp8TTdOTSvcDnm
m/zsLPE4WkPmjPIUmXuerntxnMAtnQy3hnNke2/DZKuNtZt+vhI7UIJBcYdE4pXd
skXlxKAQD/07b0cfm/kIC94gJEeiYy9DliTxBiFpQuB6NgJi0W+pmPdjWKmRMm8H
5bW1oOn04hOUOqCGk3RQM2hkHJLT+2Q/KBf1lX1v+VF6paCKycoY8FpxOIZf9xIf
0jJFv3xhJme0ldxv+ZK1QWZxRWd9dA16CSfG4JrxGj/bgZzEEbG5v9nmuwN0Ra1u
BRrh+3DLdnDMZ3gihX6AzrrEg3Sp9pj6vSMFAvYMkuXSi8VtwniGrHo7E8mNPNIG
w1/41TaiyEIzNtLMqBqibRQYkf20s07bcUjQHhiH5x/1xASnBNWvV24mJgETMjCI
Ddro6qiJjby3cf4rAIypRRx1IlSVeCZvOvnRfBOis/lWX8t5zu5q3UnlDxm2jmn0
6V4iIjBYguNjmGvf1uSRDF7pMTYSzBqLeAcGeDDk144NXL47+EZGXpOr5zKmGbTX
EbxC9AdhwTg4n2KcveSCiiF1kECrF7rpyn8A+qlaxtacxRRipx1huvvIQnP5Uxdk
dNLIqyud2+uYlbSTk4WxbNJo41UXCr5b8YR9JW98VtoZ/J1ORTWNoeXdkdcQA5NU
tjt5rSAUaksAAFWEUa+aL4Xa7XRhmA6jsBMLVp3kwMcWIAuZMMCY2xD5TW0e/lQQ
1dAmx1aItpWKMX0OWq1RK9Mh4+h4GHMhmimuLpfe63Yh7YsNTTSLUwBY/QCVtfYi
/yToMfPlXS7zPHbLKx+He8TZNiIGX4NM686lbkK1QMw77KVfTyBf6LVe0J8bA1MC
szxwSuqrLOLgkt2Q4pOROdmEsYT+3TEANFnQly6+SPQI+n4Z0YYdeJhmDYeclNrq
SgembCav06i2/FBee3GjsmzfB0CcQe/41EyismQoJuv+dK9d6iHZXK3bscEwoQIn
zSVOAkEAo+Bp7aYpUQ6gHyGASuSTpQfdcDzG4sR7+ZDK4PTOMs6R78bUUv5qoyj0
y/t96nW3u/oS9OEUPH2xjtlHkK+QhwYmMXZ2pbhWtUno73RcliAnCuiE/to7jfmS
eCgkfaqBf/h+tgMstiKXuP8RAcOip+8R/4x4DqjDd+hxyVatTCtLc0WChgjR0DWf
ORIFepzDUz+onMHw3lTfaT2oxHqg73QKC9QhnyBrw/UEXE8FI1Vjro3H9sqXZ/wl
ughioOzzisi7+eQ6C5nwf9K8ac6VNox4CP+k1HFJ4QeMdODoMgaFONOeFsKm25VA
l4AP3PlvWH/pegeyU3cpEd7XL4fFIzZgRJAG2taQTyaFsZtHJmVvK/FH6mRRFS0t
ZlKqO9Y5JJthCA0mLe3gFNDrul7k04d8HK8QxZWEw9BWA+pX1NTnjczE6n76QGk4
Y6xBN5KG2ubO/zh+1pmRM+VyBE6BoX3CU72FVjhKzNxSMx/JtpYSELweI4ArGEHa
tFr7+XXf3jT4DEECOVSMUsWtrQIkOlmMnGLwcvPUwm5SZDD6uWHvyKnrBEy+fqLG
eE2XaiNF9yvCItQMd7CakUkqBZh2hPngWzPglB0pU/rx3PG+ds3Vj8fMHcG7Ir0p
x2RKWNFWBtUhJe5ReVPNO0Z6+J2QPAf118BcmY33/ZLony8udcfwls6r+R/J2nNu
JePRk0wq65NofBYTpI763KHawErEJPMcGy65Nofwg1u5r5G+1sup/pXq/8XNFcp2
VSTAbyR7v+0ZfLBxz2pDv9M2HzTl2UiTdKyWTA+xzu7KVvGasSe3dtfAxK7flSmX
6+iDwPDaDAOpWRRm1yz5+0iSCZbFKuQ+G9QHfF+PeURF8hhPD2DKh8/UDnT/Zxfj
mCTTy7ZKx2E8VAZrN/ZBvf10TUZUB6te6Sj4igNX6XfQYWu/UkUGcIk4+4sa5RTp
cBjfWCJocpD0ma3MOdHzZc/Mkm5Q44dtJSFZTgRuIie8c28HjOq2CNhMO/ebWwpM
LM9aYWEx8EonK7ajuf460ZN2uGFBq2B8JvMyo/qUmFNMHFhexsmBkTKYFQZDXsR7
iA2Gj6gHwTc+bMemclg4U4NTRen/vppG6xSqiPMv7FieMCtbLwpVrUJCwRjHX0T3
SEMKfDq0VsPsBZbwB5+SSJvBU8z3TRw2a0mHcnAZBFU23h03Pd2QghVA5OXtFUAv
le4ZNl81wXvikFRyz1hm9EzokqnEiqUa6uZxv1ZyZj5lBV+WqehraD8DRljr1WO3
xEKoSGCTixBnV6CS3RGaqlAn4uLb5dPRyyfesiFV6WqZFhtUXoSiiR5kyrkcPaOy
j44riu8NtYbLsxcyQUcoXMzYsy+OK9LIG8RIApyKrSiV2VHvWAdvjV3mzbsrlXoP
3xotuvxvzuDBDDFA19wPmZPosHK13QMmkMUDZCrjEe/qnFCOwsMaNrVN948Ww2gA
SYFqUJqST0JZr57eM8pfhVjwju0RikOH3gMvzF7fEturC0N80vX/PeZC8lvFq/1v
wU3cc4H6YvrvwanSXWIdH+3LhpzGWCuSRpgfkmjY1hXgDkRzhupBpVK78rFDKFAn
eVmTvU6bo/qQ/Ulta3X7f1e+qC7AtkxHWim+9WZSK8+9hDSS3Rh00FXxw3qVflmj
QsvSEGrcux/UOI+XbX5nUJvuNW/qNrL39whOO1Gv79HsuyRD7EInqVKMF9P+jcRy
6s6JCldBXngUSE0bYhd6Inggg6RFDomFCyqWxddke1oJndP/PkpevNLFzXcL4sAB
77P6bVsa04VLA1UFyXPQFbjaHnkw6C48dJAeh9Snn9BtpHfkyjHJh3LUSoFbz3px
ZFjs+IQofEpepHr1PdzRBk2bY789fkBmVnoRWKHaG+x7xDrGSNzx7qRcERE2o30d
bOIs25gN2mI/myOT986oHgr9mznBNGKPEJnuCMrBJPSWfaWUYgR/+ncQYvT8phgT
JJS6YysEKQj2EYsUr0Zo1Rz5ihDhtI2AXdFmprH8ArCys2UAHgTsYJqIaB1i5J6E
KQB0bVhgDCNGC7Muhrgd7QA1KOr4SUtr6x3vdF8yI7a1/hvWkYoMMsTNbjHK+vVI
VEZtm21GheGrUrkBqBUeFrlwnJqmoavTRKNflCKlCwvOTgZ7qyEW5ev5jLX+IKCw
yxE2SlHd4JLjiC7IvAx20OCtfQt6oCgqOLEsiZ5KlPNXV2qetLq6Xbgtdw8LWht2
nsbqau1A4wKzM2nGRFLC8/oPjqMkuh21mZNj23oYs4VU0vVFVLQHpAGZtctNx68D
c14LeSgJZAhQ+oUP9mDaeSknjS1IuemFRgmgSR7qyjHAB4KiytpT7/uJyYqhrTDi
cz7xD6qrbXISGVtXikkZCuOfP42GOyiF4mCl+cVqmUw1lHZPP8hF9/m8gJ654/0d
QH3TeX7eoCwty0YdCs1o57tD6rO9tL6S0uv2V/8lu/dkchltHCG5ppqAbMzUS2eu
/YTSrJDc2AtMwuw3wF3USGwYhp6aL65TvU9JMtEsvMLJfW6kgZZZfpycPCmgPUos
xhU7/rSVn4DouB60eiEvDzq3xkZ8ui7wssey1VLZs4Dk8wNwSGTZGlJu+ZLxFUah
fQEof6b2OFx5WoXkGJT3mSRJih725ZoWn/M+ex8YIsoRMD4y7pytg6viIapVY8C0
Dy5Qd8DT+mbqEHcChrNiy9mQ0EXhX7bTr3kC63rr5yehGgADxEvwUpZ3oHHYkKl+
ghQnaw2RPeiiedC7Tf2wryl7oL6JFoQZO5sojnPT5zVi5nKkyIKnMpeLUAHbs8sY
1uyJUkKfWvXwqLwmRN3YWssKhsbpdR8R7AtbLEmUshbHgnLviPNuQ0j9RHjN+90D
z4KmtuMkOCjfvuBLTRyjI0w9lDckvG+YpvO5huFFA8jXULVwFHbo242/QQtkMD0q
904gDrAxEqVcgBCHbZ+rViHEFsXTcuetxGL8nQ2D72VMEL3pO1ZhLdhMY4UYawEY
ll0kW/A6H1vH3OoYMLNqj7WRQQ4UgGbEmOpTsNgF+d8QpHM0O5NJ+8sEAGAWzTlP
mx1yprod1xEkWjPDWX80eCbnhyi2RIFUO3MWP1HbvE/RKGYViLAKlJBkD0nSAyoL
SbP8LeHpuVirfJKsjeOMtX0vrHZs/ejklhLNaW+H9j4OTHE8OtomGkhqyptFeNwG
xVwpn0v3opJVL2sc4+loiP6zfMmPiXen52nhkBq4AeCqKq4lB/k61MGVtiM9RWeC
DNZJKP2Z9eZ9gO8njgFde6ty+PrvAHb1BGIH9lolvn6LyyGpMJqdrcjK1EGy1GuG
zHqHwIPHXRv4rg4g+fdNTcGlXvemvbk3hD8Wont4YLgW/2Em1gKy0RtTygXjqYVA
WNEuJEaR/Z/84D6gHEwhEqrafOMmznj7AM9kffEkVNldgxckcRrfV1QRo9VnX00D
tb5WP2uLrVCNqais9PFtj0KuPfS+Db8OkiwbEO24YILnhOre/RDXo1Uz/HR1e8Ch
yJZggWxpWPLyJX5WM5G+t0cgZXOnJ+WaGCt48VpieexGO/knQsh7DigRGoAVUIGy
uRTKRRvJyhIvZC0TvtH3YyzNGBQ4x6HRa3ZiZ/9+fOlPCrLL9rt5p8LgJIg5jY2k
Ce7YDvsNvn9m8QJLnC8vAoNK2km2Alg6wSnypnh+r8fqbStnqwqGiiR6v4eAXfFX
AzVPkJBObifkLcgeqT3loKg3B0XYdVI/9RDyQZkIwdhkox9NX61p7pAH0S0a+3el
dhCv9uo78W5q7dUA28DfyUeZgYBClwVb8VFa8YKCT8epYZdisJaPzWktpP10hCmv
fLyEwGVQdA5oYQvi8LA8a9D3zvi9MyBaAg1PO+9pEtxi9ZYpKF45Ex9sAVD6Nvkd
V+KYaMfWHLGd+IbfN7zQwm4qP6wappBnv+0m/BcnfmylDtT9scJ9OlFpl5vdlUQM
nvojBnEdfeePxxnHekProAFYDJsabqfTdKkVR41IL0rkzSZUdmp8k0Uu0IIy7AV3
D4XMH3110WCexo2pxJ9GdniJXHozKd0O4RxQfEmQ43OjwBJ9PXBLUnif1CEGa9IG
+A+ReKYATWg/h9X04QGEfRBMISFCG+FgVMU/VPIf8Cf5FqTrBzfL2v64pPJlU1eI
p7R8/bd+hD02sidG+MgakrrHxOv9LCuuBGpcmPleC9EYFYH4f1UDdiWW2J2otE1B
tiDdInWE4cNuaKj3MhRM0ncintFFs+wckt0Ecg/TzwTGjHVYzIq1Cb+Zw9hIhAvk
ES9QqLu/Eo/J+HGQ5oTnQvYlBjvIhGF9IB2JrK87/wXR+p+AWc0HB6Zlmvwv0fMQ
wJLkVRH745Y4lqfKRmzjhHsWfUce3pH0MBsV/lQTVCTtsHsNXSXN00SHDLaYo3wh
HsWOt5n2pgFrJc+uVjkicYkii1hdjik/s7P9ftkhucLCEjoD5xrbU+4T6cfiDzMo
XXFxZgKVoswGsCBC0DwMt/7Jx1u3BjYUC7W2amS6uchiTKGMwO350CXgJ3XFIuio
pN517zYebsyEvDUV1QM/Onv/m+eR5rXA3axn2fvwCYC0KePX6Lie045+jm7loDjP
A1/RCnvoKRyrFN/+jejhlX+DOAYkNHcQoitCYsk4IrNNm4PXaRcnL8xtjB969Zmx
+Z9/aJiFtYHgLeK/PG5+dpSZsLfANcA8PYTcbUiwdK2CgsA1/O9B9EkgU5L0tgFh
byE9G+Z7gKDvukOE758/PbwTRNGG/EEuXa+OywflX5Wfpmy1DiwTYfDeaYtxL27s
8VMj/8m51mjQus5hI7YIhngq//6leqWdWF6TlExxElMO8au7HQlqbemxol3h7J1B
jIQK7UAdE+6enRr82TwFAYxAgppvw6Ip4HLnMKNTIWYG3NfTkppDFF63DtfebWMD
UR6MvwHwuo0jqpnLFB4zvf2GGf7bDnK9KjrEAUDQ+dULKWcUwjpStGoExyHqWUbD
pBZvzQwsAilEKH6hMF2wll4DTGMoKkcgRBJN7EV2zKTfP0B8JOjtBj4NWM1bs8Ui
sG4Su/VwLAgb//XTIaXtfH9dCo9Eyt4rndGyfRe4Eutyr0BRNSYjHqfqgXYKAZGx
Zh2EVzKtU+op2zy8sfIPIn+0e2mwl6Iq1YicGxDnzMc=
`pragma protect end_protected
