-- sdi_ip_ii_rx.vhd

-- Generated using ACDS version 15.0 145

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sdi_ip_ii_rx is
	port (
		rx_dataout              : out std_logic_vector(19 downto 0);                    --              rx_dataout.export
		rx_dataout_valid        : out std_logic;                                        --        rx_dataout_valid.export
		rx_f                    : out std_logic_vector(0 downto 0);                     --                    rx_f.export
		rx_v                    : out std_logic_vector(0 downto 0);                     --                    rx_v.export
		rx_h                    : out std_logic_vector(0 downto 0);                     --                    rx_h.export
		rx_ap                   : out std_logic_vector(0 downto 0);                     --                   rx_ap.export
		rx_format               : out std_logic_vector(4 downto 0);                     --               rx_format.export
		rx_eav                  : out std_logic_vector(0 downto 0);                     --                  rx_eav.export
		rx_trs                  : out std_logic_vector(0 downto 0);                     --                  rx_trs.export
		rx_align_locked         : out std_logic;                                        --         rx_align_locked.export
		rx_trs_locked           : out std_logic_vector(0 downto 0);                     --           rx_trs_locked.export
		rx_frame_locked         : out std_logic;                                        --         rx_frame_locked.export
		rx_ln                   : out std_logic_vector(10 downto 0);                    --                   rx_ln.export
		rx_clkout               : out std_logic;                                        --               rx_clkout.clk
		rx_coreclk_is_ntsc_paln : in  std_logic                     := '0';             -- rx_coreclk_is_ntsc_paln.export
		rx_clkout_is_ntsc_paln  : out std_logic;                                        --  rx_clkout_is_ntsc_paln.export
		rx_rst_proto_out        : out std_logic;                                        --        rx_rst_proto_out.export
		rx_rst                  : in  std_logic                     := '0';             --                  rx_rst.reset
		rx_coreclk              : in  std_logic                     := '0';             --              rx_coreclk.clk
		xcvr_refclk             : in  std_logic                     := '0';             --             xcvr_refclk.clk
		sdi_rx                  : in  std_logic                     := '0';             --                  sdi_rx.export
		rx_pll_locked           : out std_logic;                                        --           rx_pll_locked.export
		reconfig_to_xcvr        : in  std_logic_vector(69 downto 0) := (others => '0'); --        reconfig_to_xcvr.reconfig_to_xcvr
		reconfig_from_xcvr      : out std_logic_vector(45 downto 0)                     --      reconfig_from_xcvr.reconfig_from_xcvr
	);
end entity sdi_ip_ii_rx;

architecture rtl of sdi_ip_ii_rx is
	component sdi_ii_0001_rx is
		generic (
			FAMILY               : string  := "STRATIX V";
			VIDEO_STANDARD       : string  := "hd";
			SD_BIT_WIDTH         : integer := 10;
			DIRECTION            : string  := "du";
			TRANSCEIVER_PROTOCOL : string  := "xcvr_proto";
			HD_FREQ              : string  := "148.5";
			XCVR_TX_PLL_SEL      : integer := 0;
			RX_INC_ERR_TOLERANCE : integer := 0;
			RX_CRC_ERROR_OUTPUT  : integer := 0;
			RX_EN_VPID_EXTRACT   : integer := 0;
			RX_EN_A2B_CONV       : integer := 0;
			RX_EN_B2A_CONV       : integer := 0;
			TX_EN_VPID_INSERT    : integer := 0;
			IS_RTL_SIM           : integer := 0
		);
		port (
			rx_dataout              : out std_logic_vector(19 downto 0);                    -- export
			rx_dataout_valid        : out std_logic;                                        -- export
			rx_f                    : out std_logic_vector(0 downto 0);                     -- export
			rx_v                    : out std_logic_vector(0 downto 0);                     -- export
			rx_h                    : out std_logic_vector(0 downto 0);                     -- export
			rx_ap                   : out std_logic_vector(0 downto 0);                     -- export
			rx_format               : out std_logic_vector(4 downto 0);                     -- export
			rx_eav                  : out std_logic_vector(0 downto 0);                     -- export
			rx_trs                  : out std_logic_vector(0 downto 0);                     -- export
			rx_align_locked         : out std_logic;                                        -- export
			rx_trs_locked           : out std_logic_vector(0 downto 0);                     -- export
			rx_frame_locked         : out std_logic;                                        -- export
			rx_ln                   : out std_logic_vector(10 downto 0);                    -- export
			rx_clkout               : out std_logic;                                        -- clk
			rx_coreclk_is_ntsc_paln : in  std_logic                     := 'X';             -- export
			rx_clkout_is_ntsc_paln  : out std_logic;                                        -- export
			rx_rst_proto_out        : out std_logic;                                        -- export
			rx_rst                  : in  std_logic                     := 'X';             -- reset
			rx_coreclk              : in  std_logic                     := 'X';             -- clk
			xcvr_refclk             : in  std_logic                     := 'X';             -- clk
			sdi_rx                  : in  std_logic                     := 'X';             -- export
			rx_pll_locked           : out std_logic;                                        -- export
			reconfig_to_xcvr        : in  std_logic_vector(69 downto 0) := (others => 'X'); -- reconfig_to_xcvr
			reconfig_from_xcvr      : out std_logic_vector(45 downto 0)                     -- reconfig_from_xcvr
		);
	end component sdi_ii_0001_rx;

begin

	-- sdi_ip_ii_rx_inst : entity sdi_ip_ii_rx.sdi_ii_0001
	sdi_ip_ii_rx_inst : component sdi_ii_0001_rx
		generic map (
			FAMILY               => "Cyclone V",
			VIDEO_STANDARD       => "hd",
			SD_BIT_WIDTH         => 10,
			DIRECTION            => "rx",
			TRANSCEIVER_PROTOCOL => "xcvr_proto",
			HD_FREQ              => "148.5",
			XCVR_TX_PLL_SEL      => 0,
			RX_INC_ERR_TOLERANCE => 0,
			RX_CRC_ERROR_OUTPUT  => 0,
			RX_EN_VPID_EXTRACT   => 0,
			RX_EN_A2B_CONV       => 0,
			RX_EN_B2A_CONV       => 0,
			TX_EN_VPID_INSERT    => 0,
			IS_RTL_SIM           => 0
		)
		port map (
			rx_dataout              => rx_dataout,              --              rx_dataout.export
			rx_dataout_valid        => rx_dataout_valid,        --        rx_dataout_valid.export
			rx_f                    => rx_f,                    --                    rx_f.export
			rx_v                    => rx_v,                    --                    rx_v.export
			rx_h                    => rx_h,                    --                    rx_h.export
			rx_ap                   => rx_ap,                   --                   rx_ap.export
			rx_format               => rx_format,               --               rx_format.export
			rx_eav                  => rx_eav,                  --                  rx_eav.export
			rx_trs                  => rx_trs,                  --                  rx_trs.export
			rx_align_locked         => rx_align_locked,         --         rx_align_locked.export
			rx_trs_locked           => rx_trs_locked,           --           rx_trs_locked.export
			rx_frame_locked         => rx_frame_locked,         --         rx_frame_locked.export
			rx_ln                   => rx_ln,                   --                   rx_ln.export
			rx_clkout               => rx_clkout,               --               rx_clkout.clk
			rx_coreclk_is_ntsc_paln => rx_coreclk_is_ntsc_paln, -- rx_coreclk_is_ntsc_paln.export
			rx_clkout_is_ntsc_paln  => rx_clkout_is_ntsc_paln,  --  rx_clkout_is_ntsc_paln.export
			rx_rst_proto_out        => rx_rst_proto_out,        --        rx_rst_proto_out.export
			rx_rst                  => rx_rst,                  --                  rx_rst.reset
			rx_coreclk              => rx_coreclk,              --              rx_coreclk.clk
			xcvr_refclk             => xcvr_refclk,             --             xcvr_refclk.clk
			sdi_rx                  => sdi_rx,                  --                  sdi_rx.export
			rx_pll_locked           => rx_pll_locked,           --           rx_pll_locked.export
			reconfig_to_xcvr        => reconfig_to_xcvr,        --        reconfig_to_xcvr.reconfig_to_xcvr
			reconfig_from_xcvr      => reconfig_from_xcvr       --      reconfig_from_xcvr.reconfig_from_xcvr
		);

end architecture rtl; -- of sdi_ip_ii_rx
