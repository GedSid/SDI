// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:37 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
e0NgIsop1sM3IdxAESSuA5iEzACJ7DI7Bt5M/jaZJlJ/VffvAHx9OxFGsGEUlYtl
TfGInm3oitFTmI2f337IG/YvNSCptapqCRZqZ8LiWWkxWL4dL+xzCPRSdyeFk07s
FOEYkc9+kRYrO9UiRwjnD4f5ovQjrcPl6pAuaX8ovM4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28224)
zinEEIN0wLncRtcYNzj6o18iVqhhxeZub4JKgvkHXE/Je+VldhsZeHwNhOjVQMFl
k5/bfhOibW4GpA49oUsRQ2PxuzriNRGIngcY5EqC1l+ulmw3KZztnm62xmkEvVWa
SUGc1WoRJyCUpLpGIOniSqfErW9wdZ98djm7fYTCPLZ6RN1F5L1mL11qHswMrjk7
lnevRkOwKO7TWJ7Esn8fz65dXuOiX5kUx+9c1hqXa92hPcfe1kKa7nZXxfpg24kU
u32bQNDIqfPFpsq7CtgNNIrVbtZbGT8v3teftxJgfr/FNrcTgePDVt8pDN+47X9T
VfEmoEFl40eWwHu6vC8s/md5sFI+fNzswNIhI65oDUss9p/VvDFJx0Z4svJjUjFw
E0OIUftUGn5YsHE7+9B/eCZsXNxeikRoZmvARlpj1dreHCUHEuyV2OVxOer/SbJC
batDon9ypKAW/Wc20uRACNvlRQ/ICHS3NZf7HLSXdgDWdSUkYaLFElP+0BZDMslN
mrqdc6pwKBVNqC4/jlHkMsAvWH9hTN8l9Fno3ZpK7huNJBOUtFuSEC/5hi7zqdlI
bNctOXekZ/o/ryUcH6AgNYcKOb0mVJamzkqSgl7OaaqQW9nZ8b/T8SCJWCV2zD06
tCLodjIgPaZFBuUMr5zu/lPwuVGX0K6gLzTeUF0KKCuL8iHGb+ztPU4dVYxldIk9
ZzgzN8OZM5n3yr5o1O3iQUQfdWlbUFt7bN82MNwlsZXFPg4EkdbtTAlrNYnD3F53
DHnUUwSCzioOHTypMvfJrIPaOoqAjLncWfsM2tNQFYR0te+3dJD+BXUklsFNLg33
mnN2IFUDrHrOt7bCNa0cWLcirXM0mQm7lyUMITvO5Zv2jQxlXG/9q5aJs/WvdBn0
YitgL9CaaOGHeNULVusSBCiOkJxxwNTk5g6T4e7UqKvaaR7iYzWv9NAeCL8bVllW
2c8X7iWQz0kgH5KREHpelIqQXSh5fvmmP6eXT/q//s7Pw/fh123pNcFe9sV6Ya9Q
+H7d/7fOoazxvDW5+7C56vKoaNK29rtJ5BtFfGcDuzmlmeqlxUG3fggVOgN5Zo/h
+quz8dmxWKXrIxrU7jW08g1sI8aJA+7N2umWzW11/+p9OLcmrcy37LY87qe3z8v2
lzynQQdj+5gp07FpsnZAyhtnLAlz0gfbWwMjhiNM0WOT4fAvR67ERQNDaH5FQUzI
RVCCeBUP9vzVAhFdd2bhmvzw/0LH7Yu4sXtNLooGw+1JbrKAJkoLavR8QNjdq29s
B2kkzkJosDvOPzGITFDLr306HpSdJ6UoCcrVB18boHJOF3TV1ip6BeWMQBLOIwuN
E9NHjmJQqrLtEn1DHeJi0m5qletLojpP0+jXwbani/Ege2/xV4U/gJXzmAV4UY97
2vviJwTsWzQ33yZAqCCtvYa7bvuyXqgA7dj65HGaZjq2UwFNu6m3JNY4yWIHgU/i
t5xSHyDLQxhko8BSfCVL5MDp7t5AQPuq96nrj7UCSQpwlpXRFdemzDGlkZKpNmoG
yANBmD8tqAteb+f0wqIjBaKo0Rj9wwop7ggupAozpjdm3uMdApypnADAqjVsQJ16
aJMHxOfAsJExD0814jLQ19sgJmLZ9gwcvg+SVA61a6du+mtLnfUnu3jFAHjXR3XB
AlbWpt9GXRSh0Nz/YCOJOa1pcQm87Q+mRBBwcXeavCqPE7tGbz11HzPP+i4CKntp
zY9T+gB9PUkLxF19b0YBPfbEdgcHc4jj4LHHYp1EEz4tiiL7EdsthxX70FAvqC5u
zSi2eoysG7nQtvNpRiAKuUjd3b+hFfFiOVn6+y1Aef0tdXomXIiLrsG5WDcqrjnl
ZpvYXP8gP50gQARbCpMomuOU+JqjmVQi0Y4IXqXtejgDLkWXkcmC0oVrCZ2Lst8p
tC84QbeaSruNr+6ppmRAg8QazwKt8ACwtdgmPzTAvRz8z6MzEOvq2AdhMbsQ6JvN
ocj5blW3WT3SFksb03NonhYQlohdclwFzm19Gm/9AOsMfnSkVvEnPCbqu89HyN+h
+5Eqa7PHhSeYfJHft44/JrebAt6efPwCpJdBbLRS5h+GzMtWmS6sCZxlJVSs91AH
VoQgc2A7YDMYoFhGkvYQxGLynfJ1zUcxLXggQxMOGPdfRO1pKbZ/r26nimyBB1D1
Tgt7EedVrQRhckqUDGiaOkoLTf7G32xFrH1IJdJJCuTWqPMnOa+ZLBoR1tbUlJVS
3ryNnNIWY4+2KcXlXzWpBC64JKnAY2pVhg8ZCiam5ZpCFtOvJ6FYGVRPwtx5RVIM
1MwVNJfhJISE9SujRpsYCkGKyx0t4CfWf2VL00y+mdinJYXgcfy6zhykq0ZAKecn
5Z7CWtvZOzl1JkeofQEK45cUmSYPfdle21g8YzXiUKnawVihfnvIgGqInnkQeKcN
nNeBhXcfBEfyIbOmawWi+RhK5jM1yTN6pf+KPE+CZVPtMSUDfOlEnO2RmHwHG4U8
j4Fzs9SBAlidTzdBTjr5Ofb6g12Mqbky5pW2ivYD4A+M8vockxREg3kJKMCC/S38
LBLtBUJ0X0TSUMVu776jI4Zfodl8KMwcFqxHe833m4wrD7h/Mskux7s1XlHeYa74
LKlgdkT//l819nRM72MCt9HoxNBW4jR7VmAnfs8DQh7HcHV9NPOZd/tDrKG8y8lH
R5cf7w5PAe+Kg80kFL7aNOyf17rhJM6DpXon10reUIGAe9PPxSEFOvYBm19A+S6m
1dVig3L6RSHxRfOjzzXPOF1PYKNX8xORyvN42tGdcTUjZCA4LIPLnRVZqAdo0xVT
rfvpPjEeOvCFnMtGkL1DYuPVxNhen2WS8vcUjCDOkoDu1ssmzlsJb5uv3gpppm0d
//7zGzjkrtIyxS3zaj65rT7S33q5PkXC+ocYz3c+EFwXA4fvNL/ZflYZGLdDk5O6
h6ljXS29baZvua+rICofYRlEhIbVFDoHBibRKoznF2a3XQ15VZ9ER6vZ25HSZgj5
dltxH7vFdvh23yctgaJ7bATauhFsAqasRfMDjbQbdfC6XvZbwruF9sjZCHjeGkbZ
X88lV4Tj0IrLCmcFlvlLpwGbELIUIVOtjypY29X6N7/0NsLQaTKXR0yQnNzcRwTe
mhyX124H+U3OcrS8oFZexvaDbzIAWsyYf1cLu0mp5R4BM+fiOKeXk+ldaYXeA18i
DOMvj669khADa8z8jjsRPcN3V7IavajanNObCW0q4fni1J/DFtOYMiKfRdJ85F36
X4CiznlsWSb4/6MHsjj01AuqDPfMSQ9BFiFofbTRF5qUHv0LRke9FIeAsG+suNv/
4RkEfnI6jtXnjQPe2IAW0SvtN9tIYcrIaWUua8i5AsvQp88AxQjOv0+EYI8ljcJd
xZDuSV8nhQXBhnFeYJByyKXMpNBnzRQemSgbIIodtgB6EKEMJTdTjLYX8RHHYsN7
7+IxrozI9I5PPekvnAw4u3Befm6WRC3ZZWZoQReG8ZE8Xf8qU0IcSw5IinRsVftI
m3QqkdIXFa6CzQePzsdzy9WBbw+rg/CkO6uoPWJ1tHqfZypfD5GpqH3XhFag3nIy
FUDzjnWZ1D3X0QOFaaM7Bfm+eA6jH+Rr0XTjX1pnHVFhMdgg+mxTy+2+3DjysiyJ
tlTiKOgrokbIzYBS7fwzlIkOk0vlkfS3RPQh8R2MU+liv8epaslHReX77GfZJUHl
DrZEfo/Uh0shYZqXo7MsP6LM2I2B7FXOiuQ1jvsYYzgQtEdouzPCbEuzgXCnfcDa
/0rfsA0Y4TpeOzmSqOhpvSqcGHqndmerk4rU2JgjyvV+RKVDzDy7JCwvLRdLOBMS
QFOEjHc9rBBU6myr8okq2YHx3GQOthSl1ype8Bc7G6uCmlwPzLyG9ufhUZg355l3
t2GkHbT/ktsX36MaCD5oa3ZiBQMLXmiBrcHnxJT0Ugzxxh2dWIKQfHtWzS8axAOh
A5xxHSgWUhiewWs5H2AxyATHGOUvP1mqg7aTlpVq3rSraj3g3z4lfNW1n3ka5e52
E2pM+4L7Lpn4mZr4P4DgldOG301DoMvrSRJbcTJdIgSL/VRqHP6f0EPnm/6+lor1
58aOp5aoCnJhqEnZHceCacMBrF+Q+pKULLPqydaM9IugNgXJJ/xFDaVnNEjgv3g2
saSg1Zao+NUyjAu5b/FVXLspPH1czRlhAbBcjZ/9PYm/y4XZ0DKDCbR6E9YEc3bO
iG3JZU/BAkmOyqfQROkpisRpz9aSZqUf7qtJAeZAq/rrpCxQPuNUeCJCz9zG4ewf
SRorDucePvbB++Rw+M+e0+npN0XDNwZiIFpKEtDpkJeRPSajFs4t0++agzs5ub9Y
zxEPSVFmBZfoVUsH25M2yOg0ZKQvs4lxi2hv7Phkmh9ZzU8d7X9720rJlQfupWdz
alHuBCRJNeaROcf8xngrFTDWDWh1fFnl0ZtsONsIcjRoiXHT/+IOC99oluQnDtuw
Ubgaj9N98WkWlwR+6byUvc8mn6sfOUZTBbJfpSm391nwWn/0ErdJMhD/Vz14P65M
X2r8mwDiMCi5rUL663DK9z7/J5MLJ7CzMeTttUCmeXGog47IkiQuR4fmfeze+E3P
pa4S1F1RkP/PH8T6nRxupMdDFsFp2bogkuvGuIc2hG9JtOIdCJMSWX9T51DYE6Ue
stkZ09tKb5qVh2K//k8DKQeYryc5WN3IilfMPKfFi2uox11+v8yA9qbaJBl5orX1
F9T4DgX7Eg/U8GNpatRtl1xblziqOgFLFtsQSxF8pQ//xFxgNA5udCpiOjzO/lWF
ghCBADiywcxwCINqkXiQtP6yKb46EjB/GcdqOgBad0dZuxqKmwQQHUVmI5xU+SJT
LMV5DvboeVut+n4q7hiTIz80aIZdzA4iuNKO4yFJk9azwXLDPxfj8lt5+MbIBiWd
gv36QpqbebQFLC2ufomLSFXH+ccKNMA8qro29xka4VaIgt3Y6Hy+Asy3Q69i8GLb
GFD2aIvfKLo/BnHRWttZkmE6yUiN1n2u9gHLo2UbRowi9oSr84xJJ+7GGjBuQ/1H
2o43/CBpAhAWmmOLPVAR2yzo0cTF2kw7hjIAHgcH9s1sHg7ajQ+mBMgBabZaDE4G
Es8TSmweiKTS2ENxiD02zIzXRAsNJjeQjNNfvqx/zdP0xtEeaKMsXuAQDKOkQRK2
rzw7JWXeEkPP/OSdMJ7J8umN56cjcy0O/+gmo8b+6dhZStbkB6blNWrb3UStDywO
CVdtUG4FNb6/0ELKH8Tp41gUp+Xf++q5Ekll7roiD7RU0hcJdDAZ/qZQFiDtAxYq
gBeE1OAVscLrfUv2CwWFQ/q8QAwFs4Z5Icy8zwiItgtFEzYaKiEx3xWbniZD6uQZ
nSFG772FlBcpPDFiGL7uTKq/L8rG48FZii/utU6qEQhfFXY5c4TT6EiYXopKsHr/
cFMqu/SlablpaIDHEexr8dfVOcv84mVHI5HZhhiq42zgdsDWGpcTzvaZMKQ5ZIsC
iLfNhd5c3cJRI2OPuS75LxwrMHkbXkJgn/IN8+J4uWtbSXuXK0tX7hqF1CUyY1VZ
g4b0m+VrHAuKuc456jxU4ZZXSb+ZEZ6m6/IhavOdC1/2Z59YC5ADXlm6mNzZLuH3
jMs/oCLwpxLYCg59cwqzjzvTcxzPfa4bnkmSI716T77IdWaGkouuiN7ozQipLFTy
t3MtNDFZSRHq4B2qRzgTId626iq8wU+vyHgkgCltbKJGMYS/CeC3dnjDm+JK8lfM
rZQdC2ksA7AIGujWdjvUikzJRjWJmUYPVr3q3kvASFUWeRuifg6XcpvSbWWnB2ci
C/HVSgtNFt0Jx7OVOl7igpI2OyECFO3zcFYx7gTvmTva3S8XNnYtBD+Vti1+CgMV
NcIpsmM+jol8d76YJF5w7vo4R3BAyyHtk7a2iM+hWGwc6y9RY9O+A7/giVZ7njpA
ESwR9dbA1iW/xnAPE3eIQkYl9chi78SqmtvXkncYpfAPnWIoQqOzDUFaBN2aiM/p
ODlnNPJmHJO3I3EF+wNAqU7dYO97MynbPwsscogDS5shAHiofTpyg9bSpMz2Rk3Y
5yf82zn5+U3b7xYbPpwTDUTAOmml8LjzhBfXcQ5g2zbovywVmq3Ly3Fj73P1o3Wv
8YSSnzdYTjYzU7LUVUJTLEBN9r4s6swRnaI0SfGMOOLdvRpIyYqndxbu4Qw0zI6x
pbiv8SLEtQiTPjEUvHoT59PEwfsshYs/dD4qczyebf5VT4hWcc5w4xucaZQLeilJ
4h5c0AY4YACzEryRwKVmLigTlf7Bi1M7TO70xJVamVUzFVbOUUFPxKpYgfRr7g9C
oMTh1NcAIhRr7DDllVMza7VVcEbETX7W+F4GTDXewzZATLKe0Uduq/uR+41AwhyC
PF+zHYgVGneTw+qMYkj1OWtM/nWeiIYJ4QwrgTxX39wUaFhBVbYwjB8wVJpo7d3S
ehx1s6Rb920TUATeA0Y6BId5qBMLWV15p4YjesW44+XO8wvu13hS5AgoJfTdSV4e
JsQBh9PcS8/1OBC2p6XC3WwnVrIqvNLrHmDU2NzILzQr/xuWwlWdgbCxdczIdkyN
WheM9rTJQH5BH8v9w2Zd+EAcazi9gw3ljH2NVQlshiMjNcDrgAxdEj0ThofIgPU7
cjDT8CAT37DWv1udB4XjkBbWoAoHczE3oY0kCFQs1xRi7yR8DtcgwTBXQpZGHSC4
K0zv1IhWBl7QzlJdWxgJf23AHKvjhu+U1ggzk6QR+jbxEJoNNvW5uqN2sDECKQ6n
eDjOzTVvpdnoCQ++VVBrroD1uRTvaM644Z5uLdgdyqOiXHCoZ9AEySd1mz4L/3if
DaJr0TBd5mLIJouxP84jS40L5v9f5QIyiuOl12TlJkL/4cFC/Xn7GXQJK3qd8bSJ
gmlmQsg63BO6fXo+CgEJhr0Yx0ZITbxiWrBQ+fdVo5oXWvbI3izFrV/LjzMPFvHD
ZcpXrS8qwtryF9TudTo64raeBefBB0p6WHm3rDUEUet/kTKrWJPpGNkiIjaCAACu
2714lGywvG+O2aaLsY+UkoWhQVz9MULcwPEt1PX7A065OB19xSl7De34gx/rU1rr
EeajIZSTfrxRr53NA6lUX10myYFroz/BEu85LuESuAqSQ0o4/6d5kdie6Kz69ORT
YFeLvhpqfz1JRekGUq8KU/XVEDrQKPXs1/W/jjeeo4V5P5VUMx5vMcNhQ+C8Bj/P
ybYeNr8iH7JAiNUcSqwb1iWXQr5AmJCkAFszl+t9GMDfMVYhWGhWR43Q+StZzSnC
J7WI3/0MtihpJ4CkbU/Z/zWs9zLweBd2mP2od1lNOz9A6sROF2LHJVXviyGevPgS
L0QOXMs+Z9tC9Q1+QTaGljwdXTSk7amik9379cQJKw7jpzMv4djaCNuaS5lR5b4/
XrQzouyiEVvECpZ6cf2l5oJk/2ImzLDXi1QAA4jXJVhB7+KwMyk/HPsWtdAFQz0e
xMSivMwpIpTDdgnOLsDYRihri2OQNLdCv9XGa7Ku+Tolowkh548/aUzv8l62Obtg
IFOTBU/5T85ilTbo/1RayGRhtxt1aehTgWmkA2YTwAx2L9HPLQq77+bNVh/zMZkD
yK82Vck8tWcAiOI1apDGTt2sM+v0n+7Cc5jmOy50WGn5hJocBZzfFqpKctwAfMWD
XGbmm267TFFN5dormkWHXg2hJ1yAl5NHfPbBjDFc01c7JfEAxkjkmOO4mPmSB7ui
/senUObijtrgH0vZJOIKzOWGarEEnQLcau3KIrG0BV2E0XzjuUjxJ08Ajs/nDmg5
nOY7MXe163Ja031EkGAhC/rusXnYxLm1e6nYgdYrHlMvo8LA95U7qYfinDqc7th6
Z5g5VkYSEBlMbdi1BdVOT/5YSOOYpzCW52HwzoDgPqP4ZMbxdftzsSKZTEbbKo9b
OEjUm+sWeu/lCwU7VhdngbjjDMTA6cQ38Y+mnoiIEBx4D7D16ZkngptbqDozdPB6
0EtTHDfbkvPc5OkR5Jsbnv455aJbScgEQ8fCdBMp8HIni00Od5fDQhkjzT1oaF4+
I7Py4KoSicGfe4bFs3AO5WKo59g7cVR5i4LxfQsMv0m9uU15hOWXE3f+95ci75KL
0JyPOrtQm9N5ROkG3UUJT0jHKWH08fRXN2X2FkqE8gHJhQmdHyYSKCe1TnferS0T
QapjUihPXV6JNCp225WtoMDxQJlToqw4g4rhTCNaodHoDlDU1q9Sacfb6YOEQL8W
65HbRSnNi6a0KLml5vSzrC1rU7L+fRa7ZUmTH2OZyL+h3YOQ9p79JJGjTFWPaElo
mJSn285NO1xVN0vSvU8b6z+LbXOsPp/xsPTcX5eXYye1CQ1QNN9be4uFcoJw5Mpv
dfEde/GjazX0/dZwnRHsw47usvCWSUrnt7zrUQpJk3EuyJz8C1w/9gT0MjC0MCuP
lJeIjk4YSuCvEDn8gQZjeTzbyU9oLyEbVZR01BhTOhBMleGwixMgnxdZFKvuwd7d
LfztM+ALlxUuhf2IHQI/MrJby8+ngCJvIq2DUoyR91NVDmPNm3LhAjCWJQGHsZyX
KAR8A13NYqttadXwvYWkgF2OR3KKVhPbkwn1OAJ+nHFEDfU+5nJ0fHidMVC9WHxi
wpc/pUV8BTYoh4lHEwy+N5LYQUcPQqiJF8EmZmr6p9sEyp3QzVjTPA8mw4ClpwMv
CxIFejJ21IMfGvwpO70qk0Vl5xjwwM2zkayJqUvEDZ9Gj7STWIPQElURJYXlgZkC
3W77JUk0T94rhiAcU0Ge0hJ7qonHohjkCkAAeNpgX7IMidIb7erpo92I6aJvGUqv
vKPglPZ3eblgl8c9uwD77pAg+mlyxBauxQZ979iXnfoPDpeSH7/kKwrYVvPtepV0
71LFch6o/9aEmRI/b64+XsLCgKzZ3XqGPtj6+jZlh2jPL8DmyX8ejVMqkegTGwY6
OYJUaOqTiORWsQ2DoauSgwT7zdCtnrTouQUHQV8zCL94Zj/wPLjrsE5Ri1wC+f6V
WQw+vnA6fXBcjnwfobb9Rhmcmozit8oKOTP+YHFapFg8/odC65ddnPj4XlQBKaoY
UisTHSIWj1JBdTNxDikGN+NP+FxFvT0QMO1OKLRTDX4/6YeB4x+SwgoPJH/ef8ZA
OycB0/7uDzSZFgjRAo4gbFJGfXMkp1hQ6spci/0DPINN7FLjBb+zrg2ieCd/BsCz
wnJ3A4bKzu2YW4TJfrI450D0eYMH1rM/iRINh/8tR5EdUCieRDew07PE/3M9diL9
tBk6QO93HjSrAtO5XRVWEXIHSirGJfwrB5YI7LW+6kFfcNjdbKqXBavc1v+040wR
VCbM1+8Hj4HaiVZ/mX4cplO+bknsXQcVjqnWdYaKWw+UZiYWW0IZ7gnPAyGjvoPP
a8RL15KC8J1Rhx4h8+tiMej7Z4fTC/WX3RSlqJ6rUZe6MFw/tS65v0IzQs0Z3IDW
kSNgngzk3hMVCS4yJ/6+3PZ0RRZkZEXE8nbP/SrF9aEEizGT6c/H5EpwMrLxJ7zm
ft0Ssv544D25ec2JjmJF6YABKyaFCGK97DgDJAenmMEZrpPTSMkaA6wu3XPYbqGO
hWKaFrVC8/yClzNeQfBRUP9aOcORp+c1cCBIL3oaRboHey0+AbGLei+0O4VJIlRq
BrTJVGph8nJL9OywH7fubmZ0l9fqMF5qNTOqzXTA40cCfvP0U4ezY6S+c49FcBjS
V3+2zCk3nT/ui37OxXNFLuadTE2K1arM9FPf6N+BFb3AKRxC7v+J4o81vELvfMgg
xDuBSq1GYvOQVWSmo+rW02UW3nChBruQ4Iy87bCVm/1ApCsxZ5mpaG3oNHjiBiN/
/JI5etPPtlONbQrXPMFEdLGdwm967I6zRxZ7u+G2zLA6JbDLoSLnjDtx6H+/4mzk
1sXqeBPw0uGpnc0rhOMSkLytz6aQcBeZc1c/BMGSaCJ7xuJhjU/x6+CUXiMgm4MW
yXDvz3JGEJma/ZkkYiJNoBZx5Vzw5Mhn6jfFMw7u3NRiHmsKzSD4DBWhjfbFixN8
16g4JiFG7oxPDw6pLu++F/A7ANepKlNGI80LHCQgj47U2ppIHOTA8pY44/DirDA8
ARp+WjY8pl6Vme6YU40hLxVZarZd0xFZe787DWX+oeKYBtF7PYot7An5LbymAvvw
voCD8/DMguWxCD5AT9Lzb1f4G1Zj9h6ER40x7JBvtLdDVhIhTqcP6GHSoUYScqhG
RUN3SPMpy/2yrW3pIc+HUqTMOWxczLzLHeo1r/osa0vq7Yz0n60oaWtKGx+WaqI+
Az+8HMqOeqZVFGp/H2ABNQ16kMx+nXj0N+DsQQVyw94UqYdYD6mpopubapMEiUbT
JJA4mYHQ/J48iXcZLF9uAn0TCimxatahloGvTu6nwjSeud1Lbw05qNyMB+RZep+t
Jf0/lEoA+N46zE4NQeQF+VTcQVgsSjRjo1I88l0ltKLY34rj5gZFRuLYinyum/lv
gVQtqkDjw3wTZifDCTTQEbC0dKOr/06iodFgH8VSbbKMt0ROwM6Em5T8iKxyknS0
0Ibai+gRl8G1TCEGruJ/Kp0xeNteu4yfzbztgku7d7TBxB8YRGj5mKIUp2tvqXu3
jBCwAZd8Gs4VLNWnElymJvzm20LIyysuoJColnW7woJVZrbC4t4HYe8Za2vfGfeA
WP3WFQC2+o57jXpmoo0RozpQBM9YyFbG1sUsR1H9CVa9/vKo0RyrZFAiPWd2FJWO
woop7k75GmFMQIFMy41Y9qnthnieIzFvnIfQ1HjPkmWhrYtCCIdEhm3kAbxTgUqG
wMYDtOcU0uX1DzykMI6Fdv7yNFt2w4Al6OTJh/ZyPKhWDV8uR3PtYdr2jNPzQhjr
3o1uXAhaa0QRkLg+ncUYht3DsANB9l3BMICEg+FlsjYPoxPrRy1CX4Xx4zhuMVUp
w/3glPn1jqBROb5OJzAonZyd0ER1CT944/oIsos/fZI4Z4TI+42Lj9+1IW/XkjVD
bPnu9HQ4pbKXobpjcbRBuiAmanCuzMB05yEJPhajlAsJNYBwH+OrPUddqtZ6mOjX
eH3bmAggDJY5/lelph45yr1Ejgsu76K26wCY795U9UG7xI+5n3V6ruzlgdhtz+Nn
KtW7Ff+KylzXi2MvhV2W5JFyEVhZFD2ChHdhBCe9loo7jPC+GE4I57bli0S0eLFS
9lZ51OHm9cb0/Gqirlz2pLYA5y7Z24p5ebZUhJVWnFKwaoIf/NOVsceBlNdhVt1e
gD+NJQzk3uppv0+ZdLJXPHU7aTLjfNIabLq8mupXzEfE+ejHvf+wU0Iq6OJU8mXd
o7NjlvkuLNQ0VPd7LTImE8b1lrp4YWX19XVqv5rC+UuFTN6oMnaiidOPF9hE3C/R
t1srkwdhDXj3W+KtIO0KsLfvT5sVjkK8FdWXXiFoTkYvxESfAbOzF8G73ogck6KZ
wDjGI8n0G7a5fCx1AxDNcW3VYrmOES4p0UaSmu9Nw6nla6Vzj9GpZO67bjL+DWEB
6yhSugnP9iaAHlAIZvIkh5tgYKFzvNJB8O/mOzezvgH2XYKwJfsL0CjCAHgMKj4P
4b0FzZ6pQWoX8Zc+IrkKnD+aAu3lG1DIe0bCMzM0QYORmn7UwY4IgD3qy2HjNUYq
34bOlzMCRYqmsKCbuwtory3Kl1QZt6gJziHDCFc8shN7Q0qVg5Fq6Olc+in1SCWm
5bat0vA8e/GtBtwry2WvxdzNbgvfneMDdBT1osAP2aXJTyAknRI1TSR2Hiigrwjl
69BiO+qzJqaZju1kZ/WHAjt+VodE8xs5mSNwYoalcnXyvwMBPPJP2HqyUg3LWq9L
nI2Um2w2fon4VAE2ZZj064SAOwGt0d8DFrrAwMwKxj8dZhUsVN1IMGQI7aC3l10h
x8Z0F+NeEs8iF6zQFmGjn6QWZc/v98AzlhImIgddej33jTQsHQ7b+1Tq20FWV+xr
oMf77zBMixyUQkfcsRDZSODx8PMkGXFUAa59vh77rnbvabcEEgISoSl+5laOqafh
oDCKRtOZqk+ZL0HkTCLPHcrb383FCmXP2O8wnEJXv6eg/S9Ah0tcGfH6bZL/Ik9y
KN0WHCs/7fV5u7bEDw1lKl6nu2Z1HWhCoNptJ3DCDcvAnH/6GAS/RqLhqjTmmtBl
spv3V72ChBvCpH51OfVLZ7/UrT5o3OVTZ2YJmTRVgCsuLUiehq3O23wMoPi6LiJX
BHcQSfqqu1RnQSxAepvr9ZCsTnGC33OZun32Fvzi1q3u6pBaW/wL0R0QidSXza16
jA4xSTul5ZKT36qI+X+xoEt422eHYmbWApHLFq+ZuLBbG3lRci9Ibp61HTLwXGnl
E1wbrnFa01ug9Q8etbFOAvHJC5y68rxuOy2DzQ4lu6kIaEG1U0+A4IUPafMAG8nt
FUKtfuPb7RjF2e/TKYi7QpvIRl9helqHBzHTEuAXRnsb+8uv1DmnIDc3g/hnxVMA
xt2PQJ4J5UbIFeAtr/y1chF3aplFKvdA+ZKjJu45pLRmQkhtUYhRrPAZ5JrdzL7+
5BPhG5TzY5u8bTWT46DP0aW0kARx/U2IoiASEzrWMWrn+8dgBdWaH8LHVOx9sJ0Y
LI4usR71KWIcxqD5vL1LNbVyL9ov80zpZpxIDNUZWTIbi/NF/3DJ61TwXS9+B25f
3EreK+wPqvHOSuEGAHSneXvXh+x4uYjy9yXyJ+ztO0GECNuItwsPuFCVmif5xjjo
9pkN13ujKoF5JXTiNRTieozm0U08oV59r+D9/gfwhQw/UsFtATUQtZYu+P19NdqN
AUajGAjUUiHsHD/pjMW4c3P8CH5uqsI7ptDl2Jyfn1UoSCLkQSDZeLScgbQDcIIj
Yif9NGQSDffh/2hq4T9rINxHm+11mWj5vMZ980r3PV9/p1XP7DgVGlNNsoL+Xf/e
OTxk68Uouf/M3dxKWTXzo1XZI4SL7eV3NSrU6trwahvOWRym0znWYHJ2ZJ7l/zw5
0qu0Sqq/y7IctsFV754hFfeThtzBPG/rE9QqzRC6il8iXJoknQ+C5X1GhzgKM5xI
/Yyidhp+7FZhATXleCtJC+2TiDzXgg02x9PL0FTRWqllOKXDVOKKtijx4PvcZcp6
WIt7iIfAIirig+ENL5v25fDrMcnuqkybwMekVVm7UuNC8ycRLIeY1o+YBp+/VAaf
oYjBQyF5ZiFWBiTVvuyzAdK/pVAbUTmkVEA9NPEJBw+ayd/DITCf2EL0bLGf/GWZ
yedc7pRtETf5prpKY6aovy6kT+N0BlR7WAvD+oouSQLOJCgs7j/IrVbtC0bvMj6T
GRkj/llK+e8lMfQUzsvPUO9Y/AaGDhiFVlpZKGHaHxcSYEBzdIWRse7WW+Q/t9lr
4T9OOMScPEKCOGwvT7uB3xJQ5l8iBR+WlUTVd62aq43lxB28mJ6TCA/kH+IT0eEE
GE6bCP+Nu36GlsYvoUMkzDqfYtp0+vJSZ2Qxqd22547Uvs+UBsNFhPMKdc7Cr1Lo
tyWymOuOI27R+kf2M/EgEdVFXXIVnE30xue3Jcx1s5Eryxom2L86LDqISCIK22gY
qR2ldUbJyB779nVMzxMzaFQ0O2gJPkPSfguDdZRt5EiA8wYGB9ZwLkqKmyKSf0Iy
zb6l5t306i5Uk0CPk0fo1bsMeWVxYfhx8yPGyiiNJF4ax5uD9KHtBbypEmDkAGHt
r0oouIjiwgqAa8lkrcXmJBDnLYrEkWkJkQ+vdPFWHlw/1902JeK1Whvnyx7zHmxr
fqd8iwZA1gV2DMJSfzUPSTJ36NYyGtjLJiKv3xHT+HdLpno3M2uQLJZJFWVssKc0
dNsaq9ZndpYD8Can4d/QGs+NstNcoEFA9hWYasa/IrHdFkv/2lBqMpJF640gEjpD
D5U0xH/zhBrIeniDR5xrvH9RKQKLAWH84kpcOdREw6lE6tTrQ7oWLWYOb0L2VWv/
RuiVd1lULMfoPQdgYC9+rZegSpEd/O5EOtKnJ/QThBUxiYLcNYZ6W6CxbNgQcSY/
SCf/h9RS/6rkYxZWl48xPb7TUP++d23kWVhbQRWvF6lAP/NJUFGABKgc2riRen74
5fDSNSG5EzJBCrmWkFugTAfegxeSEMdVCyIfFzw4iOa/x+vhkGkdqEFwjtPmqgQa
i5HXmd8zAmZW4ctHgP/SgNUbPB7TbWSWBog7uBWF19VHs7lSfF1sl77A57AhouGM
VJ6MqNum04tBdsZYoJV8ffjS/H7RPnjn6ce3IF/+Z0M4zlm+fQNzibEZFyeKyUas
tgwJCwjDjv4X5pRQHFBzuFAN08rc4+MstO0VhjU0BYa1wlZ9UFwatbc8tVbbl8v+
ZlDs3LZ/V78U8VHW1acZHDJQufDL7E/gxp+TmEAdO3athHTlOC5eNtfFI7awsdvR
Vz3fyXKxrDbKsFPt9EVlLiALX9X4kO21qN9KssFsGD76GgFB5/vxz91ea9oiJTS3
bkf7Ahb53ino7wZ76lvtSe+AOSjZqBrSlWVpbjPYjixWuSxPk7fg1Bl5LvXGRRKU
X+SUzHxFtrWMAG6VZqj8u1lmVWvhzx0fUAalUbftR0t/JNjWqMkgjgZvZTZC15K7
qiN0P8rZKtLhmvlbOSbRMpICHAn2vWKRb5vWRZdBfohOX0NtObqyhGipEnfKt9Tp
wTqPcbNqCVeWKtRw0gwLJD+7GJdrZmQUaSHPeQgqc9PhhbXAXcQzzWAxwl3xPu8S
IOBtw4+4iKhh/p2JjY6WiOSk2+THcrKSo6Y7R/3i9xFpYYnp1dGg51asEDN6ZwWE
brnjguI2i1/JGEJdWouXjLXU1RaoBgAmziESw+0/6Xk78nyuQNPcLGlm+HgVyQMX
fby2IvkenQtTLVwGkoF+rM5I6tVMJhRInQK+/b39XS2oQPdfkfitxnbHUJFWcrcX
1alpqTzDRMbVkxlgbKHSN69NmmP1poGB7pkMS1I+RO0H2BROmUI2AiSMhrAW7fyf
IQ9SfmdYUbo/SvIbCEo9pzCMgCLIY2yvQ848v2XDAn267OAZHAd7unVlf+2hr/eQ
bc5T9AgOQY+sPoRtS19Hsg5+fqEHBqZl+PbixQANCrFtuba2Sfv6fV86IvEZ6AyK
9CLnh/lpM8YXnsU2E+NXuVKewfKbNGo1hJSHu56sFdDtKNqPbpigWJiaYfF6hxo5
oVCrT7SBdOLcU5af414ImeRm2Zietr6CVrJoidHrzgLUdoWb/Y8sE7qebqevjiKV
RhCvabvH6OsO1K++MFVYvDfYO0iSnjVUk3gVuasuyhc+Cb8nJXxnQ7FEMwaLkMhW
1S3w7vFZvfVzT6XsPPkkMyqYnybKorIjmqfv3tWdST2jA1xne6jtsIbpxG7057UG
KNhDkKs0+yt1ZFLkbtkaWGSkMfizpwvrbQ9TjFgVjbnO3rB05dCzQsDfahTxHo2C
QkNjplWxEJxV5JRh0L9GOaqiB8GY5ZOoFn4LSlxRgZl2HZh3FsYX4mDvjgYWQuMl
hckAyyypduknKJGryAmDELrF5elByp6ygzik3hvnb6fJ7CusVraLKaqVuYuQYz19
1DJlDXCvRfl4joT6zvRf36Nwj5q/3Dgf4efN1XdjxO0hY0n/sm/b+/r+HViorKU3
apBj90BNxAR1oJpW1DTc7qoDKbn5S/ZBXbjGMhl6QF5vfJjQA49ekeQu08aEEN5H
5b8CANy/wm2zBV3msRvhIsSdjQaNa8CH+BMGucwXot048wGRQf/dNM03B4cDstYH
SrFd4flNc4uA1Pb2wIpjUBa5oQL1aajlfgB8eaz2HBwaD3R425pTH4ds12hME+S8
P/hM4CLxBf27JsO8Ow9wgWy3ErR6bNIdWRcPoWukQeFNj9nbDO80HeC9WMkUq+oz
j1SWSKb4+4ctke4NF0ZgQF5rEO12B1Lphul/cuQSyGQrJr/kFVESRHaxjhUiAM4m
iqZASee8ElNpr4Yh2AQmPcjJgm9ljw2Ixg53FOv4XUyRf2s+H3oal0gkPhOkGOtY
DECBFBdR5wkhvW63WlwwJx0MN3IcBJKug64LEMUcpKC0FrtY4WoK35qxo/ZeI5LB
EHoJyfA/17MYzm2TvdkVjirsOu2ZB9fnR3B21izKHJR4D5n7L0vOXQ0ZdzTSWWGH
iCf6tbxicyLHGNLdCnDX/PEMK0FnYKBz/OHSKXqIyE9Xx+0gh5gCt0WEAHApHilV
qSzyrWHQvbuRsnnBqNo4Yy9Vhm+5lJ8vFD90XVFWjs5EA+IcGty+j39DrAoWrbSg
KxV54P6Og+PWHxKgzlPRdrndQDmAEFTBTg+QW0STwM/t0/Xji9gNiKUDvprUN7gE
JxFIw0po94Ke6EB5x4Vz6aUGRBqYNR+3P6/O5mMdwptfewNE7yhyj6SKEIMk9Hv1
vVdJfcwziok6xhYMAshafCapZohS2vNzH0p274D6nSY/jDGH1KcWrC1xL5UHuj9O
kOrg1wZgU2eDxaPJm2En4ncI0xt6xLm+mbjbZCKYwPXL6IHbVV5a08amBMGGK0nZ
S81kx0yJS9rFpDLYTSrQUyTSlYTIi43Npy4UspggPg1qPwGYZkizHxEqFT2JZvRY
3oK7SlEWB9tMBPP17/7Zvwyf3G/jJq1HktTxevjnSKlD9ukTe9EYVJwqB3x1W4hU
Pmll2D6vhiz26JTBl87hpgl12IER85rsbd6pGhcYb/Awt7o95Tml4SvniA5EMcbG
SRSiRtR2hklPGhTdKtLYghiFXr/udu/f3c8SKrCn5gIHMQ4bhtWIKC45SN5y9HH5
u7AUDrUSUhvnzZe1jrHhW63eWH1KZc/208UAom2C9zw5UT9n+KVfO5/RmBOBJS30
HhbNVnX8fH+VlBtrKj2mMkpCMC21tUE3seM6ZV9RmjjKwUTkGlEu2DTNABdQN049
XD4l/CTimXCQm6z6V5L5ih3xzLYXQk41harZxmv4HI7bGDKp4MVs2wtmb+hwwlF4
40XIy5lWGDGbrd5+7YY8VyRKwHHbE6NS7G7m97OcJ8aoKyVhSWgMdy6GM/qRGw01
Xx7QAclwHxX+BihvXkj91pFRtdRWbpzomoIEc+YYoQaLTyHX8Ib8l1VRN5aW+rcM
4ILCMMIC1dw0q61FSIveoHvzaDUR7XDB8yI2aEFFUCMpch5W2SgsYbUk+SzAaH5L
Q/Dfw2ApT5GJaAPDT65K2ycvB88phV2Y/DKTOm++qBIipoDI1M72fqwPvBDN+gCK
fFb6MOYYsz/FMdVrv4b4BAm8GeMFdW6E2F8ua8I27wcDoWu/kR/Vcrz8iujQfJHz
Xlyq6QW938WTUIDMWJp9RnQ9ajgf3R8q8RdKbm37HB4iVwLE+90hrkxdaFPGJ/h0
wYiNIe/qMjdOXZrVg4afBhtyT5TV58RS3Ip/ZUJA8m+9gOW5eFJX115vq/M6Ih/m
POTBD/ysjhc1MTM5Pgu2uW6T25tdHFt7RIMC3EBqD/IlWjlRGmfS+g08Nxem6fLR
a7JYf90TPAtUgMlfzOnYd2p1BBQnfOKB1iD7bBf5nP8en+cYm0NBYjmx/N+UmF+Y
xbdWU5rjWULXD69nNUeWtcPbBfqlNtRwGmLqXv4h7/bkeE1+spWDmH0rcrvr/f7F
j8G42Q1d8tX9o6LTwg/CdCgA9ykbA/Rhb3LQXZttWxEeFtTofhRBF6hFNRaPQH13
JSKFe4/TRRNlk92fdtSQXTgaXU8Wlutnf0YzZuPJPiZJyosHy629rXuhwHH19OF1
AyAMIVtNUOAp2fjGM1eptb88vBTQnzewzkGGz0vjV2e1Kyq+wq7F9uOWvrEA2RpE
3g3VCr1rL/knIyXR9dmweNtYBZDnX79gcNG0fCW9/G1eKkcGHoQOPjw58mMP+bCB
zD1muCNNfPUvCq0FyttzQnaU8rH/uZffsHfkVWsQYINddx86f3N1ECZu9i7OozFu
egC52dlHmfBvQiC4a+i3qgQgwCuDAvff3QWnT/SdaUQGigdZNu56sG6Tu5upoZT5
nQ8qVyLZ9syf+9oETQ/WAC7fo2k2/T+MLk5djMfuELGVNdf2ayjTY9slQqTSAuYu
TLxq1dvsWVdx4crCesgYAblV7/iVM382RMMkpGLU3Xv8vQ4Oz1xp9uotWGQEb0Ee
7FvU5tsXaL33+3ZDtn1SP+HgVcfqtEvMdce/PTVYx2fRVcFEVjvHH+kd12N45X50
Lz+UTlXr0vW9hc0ZB/b3AbAAmk7roZDMOeu1Jml1Dan+aOFqW5YEkGhdTco/pUAT
MNhSiIIMfTFO+Tf+wCkAO5q+rN0xkA5x9IRFDtj6c7uGOkNBXMMZzettY43NZx1w
qBeiL527/cTnuxigH+f5peNe+vBHwE/8Idv6Tmv6ZjOQNhFlIxNpBjY+FIdfCStS
y50kbkAduXB8bEqJ6D1FtWHQ3sCVuL00UmUAAnIsn6ommn2j16VmLniCI9D8Ro+K
csGO9AB52ogJd04Rp0i8wBvl6846aJMRFK8uqTjDN30xveGq4gQSbmv4RXRj7G0g
MrHbZl/Ot1B+iy0KpNpGZSJQEgg2trHza+QRm734CHzMfmVc9plvs07YlA00iphv
1fZzWvaGLj4xIcJdln1bofWXPB3jDhCIyY/JWpYzkGOSciYYFQ4Doz23hX/TflMZ
sbrfKGSMlmr6+w8awzcfpYuurahJRBFFNhVlhQqxdQ7llB8rjDWGXbtfL4ciDFlR
fE/d0nNKqNPBmkF6/x+DmPyyphYl35RXdOKp0ruL7Tv5fIpsxp9tZsq9pEiA/37b
lBDWUQLckqeZU+9X1YQmrP9dPWnpfwgdsnF///lV+XOZMhwghoM/cT6aa6cK6rgu
ARL7i2Sva3aW9yyR+dhlyzHwmTihlOjlc7LLnNlbLy7SvlNEjHNcU4i4FRzwQ025
05u852JOP5N5RVDzmyQrdSe39Q/3Gu+KTocjKNeA4nJhUuE0DW6Mn93WBDFylbcY
DDXHBfSoLEQJLDru6oDfxtJObML2R/Nj+bO0kd/PLIegJSsPK5cc4JLWCM10+/uj
8Hw2PEaXXx1WVP7hci9eIEvYoV3sXNsOEoGn2yH2SvypDtB9yOPueUzWJqFeK9MZ
Ox5N60tzWVfgFbcX/MK0z7+usbnY4YDq1on6Hh+EzqdUM/6MloU0NvtMQQff9q8S
1QYfXN6NP03PmfOgpOl4ulYh9kAsHSPwzUC/SbB6YuYt5XzrFWJKGQAcBGdgN5B6
4Cc/4qgoVXbbDanV58pkWcjp1JFXTC3W1sfjFh3B+zjPj1d+N6ff0wn7yJ5ZkpVs
yQWTpT/m15IwD/WaMhIeO8rDSHsq2Mo3Om8t+QEpOrkVjm3lJp4daPfnJ8MIBUSr
do7VeEYo1SjTLlfg1o+uXUznScQdF/+/j7aTniuieCJNlMThj0QiJHjqLIt2jZM9
b9Tc/famlKyOrRJpafLh3GTbdZRUh87/vbJogGr5kcbHmbLZrwcHz9ky7eKOPAOM
A8VZMZIpg17D7Lp5HwTJRrMFjkSMByLFyJlSLa994OhDl22aRCZ6JqfBr5NFGW3b
MaDm7N/yeNlHSod2xrTURPNLqt1u6HskXkkNQKVvwYKeNmuGN9m/GtLLTCajaIUK
ZKPDM0883TkSvEhUFtrjV+/z8ofL9xgeC986zbiC3SY837U9oQqZJ/og5ZpfgC9H
qiZhTDgMHa8NP9NtHAnkVrZ7/JLS7XzlRwjtkLckC6sHDfREYWCxWCVLg/0qxEPn
fjjjPs7kkQ1EKtEsPJMRCqqGw+XiC/JZYY3khwEH+0U5MKQWFfhjQ2lYNMrkVGmH
tUtRubKoZV3m02HEsoVavQMoARocCMu1D7BlFazBsZJa8WNcG/dwLprZqh9nfECz
EAUtwcX2J4Nma9PM5vwmUM96XYA0qRu7iMcO6EtCeEJTmb8APL91WnHq3m0d4vka
BUo7CPnCYb4zT7KMC53azFa5sO5jdJhJzoGe5dFD/GGaqsAs7SUQEYNsaElFLRjJ
OdkNuZt+RMjyjJDFVfWjL2AlHKMIxpeU9gqiWvDmGgxRAMeagx0WYsBkrRjK2SCh
Jt2Nh1VCRJa2eRamQ04QtvNKbQrEhG4TCZJroTuw0TdLZXF7JU4CqVvSHGzLfsRY
X4cdncTsQzkqBzfnpiUZcWWelp3U3WzINRszzMRMaziJ9nEtp7pFoM0MJTUr3W+8
OkmV2GKI92MX5ao10ll4hId1QFz2AEnKHqpYKiEX41veHNC6OKHtbgjm84mkkprD
oVZ6ROG9394SVQD7Mi3Cof0SyoO9FEwoeM+532B/HQk8JmZGFWpP9xBq+3bc1+C6
5rTgrnilitREiLOnU+gNH641H2SE/PbflFLxFy+8UB316gewb9Jw7aHiXWDDQ34g
sEY/nbzjo84WO2pI6/sAbz2v2Ko/58IklT7XebQhR5wTvH0Cup3vcZpAHhB7w7Kc
8BtGRkTAZkHj90Q3WGayWf/oBkAANC4NkoO7U6nacRIcl9yPe+rmUot7mzHE751U
GRAZJxRHdXq7nW0YQnWf+i4A/0C7N0qUIh7FZdwyqshbDKzOIxndiW0clfh47Sn6
18sPL6MikrJyFC3Eq5tr4LwpaPImGbBSBor4bXTxhhw9nxf0Defe6ZvnvdPWktWM
sT4i1fVjzEhFZ0oJpA0BMkw3VvBiofJfWTVPn8PUD71pp/0gOkzeht8SyShIGGH/
iwNRdVDs+SDdG1Fvo7FMvguRgzOVbRA9EjIXdiJ6I6UJQ8Ivnk/myok4tFXn2MDr
UyT38IwFue33Y+PIeyJOCLRND9MQcpShW6D30+fB+QDbbQ5MYoBpi9qJuBe1Oe23
1ex5alk+pRRrOBcFC4g8VmaY+mNmoxzraU25+cjsFszTFOpw11P9QnYKlNe2p6pU
XV6xPzsLEZohnAXMVnok2wxnzQVboeCbjqMu2l+otwn8sFofoxtFfGiWaYgE7eOx
uYX13vQDMgXeaH2M2QSXUA/uGDan09c9q+/Prbxbqe+N38euFh56OFtr9bzFOkfz
rxDpI8V8hx2ae2GyG/+JbAPN3r7tPWSDBqazd0IvrHv3C3qDpkLOP+DhpKVjWaMv
gEbgAjrrVQiit3CyYKqChk3dFY7gc6O4LTABzC+6J2PqX8OtB9294ZRekJWm9Aqx
YmsOJYKBy/kieV4OtW9SV/3o0EohkRQVhDWVURwzt8GIPOR6IzAOa4syBgpQPk3J
C6mkzJ3pgzyXII1QweqO7OF8rZJZFiaaXXBjNf4c6nVDVzoCfAAzkvriIrOGBHZf
RIGk1bu/IcLe9i3v95rmGwFNEhFXep4DNivXh1R613lkvwxCg4s7O3nx9iaacl8F
9Vag/phdt+4ss2A0fxTK1o0mEfQ3XIqFciBVp+Hn4Bcs4jcxPgln2/l9+CRiyxPk
Gj1cYfnKHnvf8brEKgj1J88fU5hWQ9yuETDGOSufEKV8rvjReFw+LAvQWXEvH/U4
JuP3mPdBba3sjz1wGFEAY8saMwsTFGieLWbNV3UvqxFLOLv5+d1XrrY6KxZW+f+9
coc51cfsWfQpjdlFulJ8F4dObqfDBVon+uuzdm49kQkN2qd3i9oQzVC3RfivQmID
65MRCpAy/KvZsUNPrRl6xpYC3/DUv3qcOF1rax0VpD5Wg5FKZRXij1hn+wzVsDZw
usSS41Ff/437oAZhZTZaBaIpC3J89b9M3XcGtTFvV2wkMfTzgxel51UMBxIvAOND
cnmh9oq0g9rEEtuvmyzrGRwOg0KjRTKnOuvxXzxr/dOyH03n8IUkoUo22WhE1kav
+sAuiQK8Z2UcqO/vHNOT6r7qHprw218gG7gXmEsZZTIFgrw5EHn1DDDj66CCx4Sg
mVXFQEK0uNl+KmJaaZqNR4meeNbySSUtnmL+vBVPBqIiuq5/TbfDdUwjkH0XWPoP
XxjrgpkLAQ6N3FHAWGJc+zJFv4qK3cs1y7AfVk+E/qsTbMv7JvIEnK37vq21qiFr
Ekai+Aab0JJTuiAlmQRl29QA7G2lA0l4KqYtWGZ1E9ksPUoXW7pz/tRQz85x3o3h
izPpRM6tm4DTrgllJZ9cdaoDtHHQ/vn8pTWfoH+81wRDItaD2YwbHXw4PD+3KfBf
ncxucqh4iWvZlBiI5mYsxjSkauRFC6TvG/Bc1lk3LBx1PJNHf5zf3UVMsGEVg598
T5Z4PdOT8cwxC85ck7hrhmB3zbaLxG5AKHt4HC4g/B1+DumFWWhS4Gk8Qk7treyX
nNlVJROVPRtBkZJoAdCLEAxg4e9nhXcmFRJ/uxNczHqljUULw2Q7A/CO3vY4uY/+
WDovx6YfKsDJ8r3UbfceEVUEUatDdIdJK1yscoGCn2fwnLuHJ5HbwPWBd4BTLRtr
vw/j9o0Ennd8Rw4uHvQZ2kPK0KdAoAcDapvmXwUsOvi64Vka9Ucjs2MyVdv/vVqf
U5QRSGCtBX18DUuKJfxHzY6TnK8MbfGUzBuBkcu54AeZr5sAHOF/Rbhas5bez8C6
ikCry20tx8866JALwmXDGK2RvOVtoHcUFQd4PeEjXbtS811wFuXfxHNM73mJq8bn
lyn/4z/7fkEM0dBQOLSVoNSjOQF5L2o0AD1641CDRz3XnkeauB2UIGjOgOnimj4Z
sm8LWfhl7iBbc1LUtd3UtZNmALsQnTKQRmosOfgML+b9ChHaS1b5jRQ8Ytq3RjJE
xxsN+xsb++NgYJYgN+0uoBs2rYkfCy+wsHnXQf62gGMWPtd56+TbmiHVOikzfRWw
p0T5DYQh5Omj7kzgsuFLOqkbfizKHyxiRmVBJA+GYrQ89ZAm/VvF7ijyu3MfuijC
cTJEGze6cnQzCPuNT7bxBqAhclibuOQdm7jBNisun6j/5e5RcDa6iVH4LwkBVD95
9RcE9yACA3MNcmtWCnSFDqYiqNDk+M7WFhpdovJH6TK7DiUCDRxx3MoBE9cEiBK6
lYslOX8JnbwKzU06eHjS6Ayn+a7CxlX6vCUFFXkW4G1nAtmfBgKw4UI4juX2TbyQ
SDkzB7cvwSHMIicskFLneTETobbZmWjUo85XHxsxD0g+eTF5OWzvV3qsmLLcPXlu
k1cAESFNb2O0kz4l27GDMgGpCUdHE04PwtOXURx8nnBLTMOfEFRjFp/5XTH85l5R
sTD6qt9OP2Nyfxndmc4Fph0TL2JIE0+52RQ6yqOiTgQQyrdC3G8r1bwGPIpVEb6B
ThkSyJicT/O6MzPIggw4eLL/UMWnJq8gy8Jaj8JF0KGCiEWoRhKbauVjthgaXZSq
RueV9xmpWIwfBbKLuTky607dXRGdoYmFXNkUigiDH3BFm/4jhIyQYNn+lfjkW0X/
eo6axjqTsUHCuwSUh8c1kTuVhRu9Ivc2ScfIv+rLXaYYyABCB+08sVDGZfu6PBXB
G/vutJsR3c6444jvggv6PG+bjLz7UPoWPrppyP8L/x2++shHw5OjcQFYLhijP0gG
AHC/WEn3aD6Jxq2U/xzUD8FgiSa8mC3hjy1fDxen/dKPYoZbrGomXFsQkC0W4JE3
1IWUPhascogFdIeoEhGBbVgT7RsyK+T5B3Me/KgcSnmIoLOrOcRMqKsPj0HNihsM
KH6f7oP0Q9LLLa95/aeYRrCVOKN6YO7jJId4vSzo1V0aGIZMyYVrVU/PrSYyXqXM
jyk6Cp6qePnK5GKEGMbaXJBBVWVVNAzngqrzW2gRxysP2PkikNO8omBjePpMOkcb
4HduS6nAH96dBkRm1t5bd6+seLeQERlwh0dIC/P2bNhoIymjch0aD5Ptmglh6jCx
MMdmvmmX4mA/aXldVzlBWewbUdgTXaGHUQAyE5v16tQ1OyTHF0jxB72NkyWI5tKM
2HOOT3eVrUG27r0TvzYH/pBvgzmiOOJLa0eRmjY2ZbPqqHm1K5pf0bDwCN3gUN3p
fdw4g3mfY8HBBli4PFny5b8qcVl4PV0vxuC50y/M94+PTEDpLa4Uox8Zds8TbYPt
VB0y/rtcw6loe4cxgDqVWmsmn+3f6L3xb15rvDSjg9TFw/cQz74dy/7f8IIBTY2d
lvIak5pbDE248xI/qF1FPLsWuGawYVoeVavQEaXuIcQPZJFBU3GkUln2iwHjmGcm
tjDHd3Bn1GTIdcpgJ/YDUv6pXOvlGL8aI+/NECdO3LyWfC57DdlWEPjpZi7bnwi7
/iC3yD8SmE6p537MJwf4QZnTYyd4n2wVVhWmVOQWqTGTSY9XuV08Jqlnle84L9B0
F8lftgm4SMQivNgmGdDtcNuMlhm9+FV7aQT/1rDawUVFpXc4XMF7k5LROiwpJqf8
7/bloan06p3mKc23M+4MjsJsqzwEVoz8gI8Mui4eT6r1A/hBb3hiRV2StplvSLFT
uxICPFCHSSm5WRHzDnZc5cWhv3sUYWA5PutA40qW4yzsC55Nd/w+4ecp5DE9DgVk
UMOu6Bz/+fQ66yObT6+Vqd6aleUOwKvS7PaIEe8+1hv6qNIKF78yFrsKNHIT30wo
Gw2T+4f78Rd3TGT+TmeE+S3piffXvJ/3h+iYWnL6KpUDSQCVBTMmF5Yx/WdCXKdM
NEQCBOeroCSc+z94rFh739OvKtPkeGHR4/MvUlmypehqjpVnfK42RnVXUGakB2ab
vfWiWhqkE3QiTMVuq5Xu7BCU3RhY6pbLcUeuA5xcy9+KgJHY+9OWvZ94dQ5jz6W2
9+3b9jOdXiUEJYyVIn/dB53XmJoV36V8djM3bgUFGGIfRTI7Yl3BnIExRkqlo1iW
eppx5knlblJ8hrMDPX8gqFpY19t7S2Id5dJlID9HPZlUuEP2KaLuewshgK/luTU3
0eZyWkfMEi8Tk2DDT79s0AnSP0Gu1ilAnO9dF5cK1xVcL3vaxZLMGTZZbPAOscpb
gd8+u3v+mv6pCRcciGTs33mFG4hvzMx2eHJq1S12AcnU4TN8raLGBbZ7LSUgIIAC
mbmt6qy2ITzmAjDaMb607Q5m9hXatOMDI2wUCLLBsPV7BWCtAb6d+YpXBlRnWDJQ
aseIq7LFFF62ytk9h/TMkRXNsiBV2lKKtUH2JxFLQKBNEswXgrQe3PIlPixWv8N/
d906DrLjjCAPfvJc6ueRw7UD1GfYRy8Tsn/Gf9mt8nniU60G+d/0RLF7JoEt6Bjn
4LRuJwV2mnx7oEMLXGpBDWvXqHarIZe9JUenqso6T7f/uFjmyIDVi5WEgzEcuo4V
H08k5sjFwWG4OnRM3FhhxVioU4NicvI4My2oWfzW8zdw4WBQoURwuLiYaXkPbPeV
z8928fTQXKir5ndMDL/xI+KSOGVMABzPrZF4bwbd/5apaCf1OCas4MoY8F3QJmkl
MKbGeqF1de5rgi/CxcEVoTaKpNltEB50fqMuFWhdj/nkaW9aZs6p+sULJv4NTZzV
C2jx10dVjWI6OBC4gzPOU85SeTHMsacsWSmRnW51m7QJvfgQITs86u525bKooBCg
x25i6K2pXTJjfjL1RIim3CBR8wAosi1uQeUNeZoQj3r+IUDRvwrolt2BDvW/B2uj
18mi2E2i12LQpSBcEPK8QCuqebb7vnzgnoS01gLEbBbMvPPuF80Fw8johvb6LB+W
mAIA42QYABSxnH3FVw/7Z41nQAADKE4lVT1WczVlQx7jWHJP8GJhssRON8PFjrP6
1S+LhqCMPzwqzqEtdxKGZXDaV3jLatMZvjZXnLFz0ZKGwjqlQ7hvNgKgOV2H+n4C
L66JkP27KQ6FBkbHbkwXS6lI4OBe5YrBDU5NczGIl/dH/dIF5W5C38IXFN28flqE
5gMFXXA+UfguKab5RzgWcEki+ciGlIR28/f+tRVqgbQ/4L9Pc/i7QaslSj8b/wr3
ClQPQ/BCUK/+1toukq6Sh1LP9KINmwHWwgcetvtyeJuer/n2VcfxQlBMgzyid1vS
cwUIOh9FfUV6jrJbYPZ6dLp+rDiDI81Bc8rOEpSo3KtWEnM0IyX9emDDCw2RCJP3
NZEgmZT+qJPQfYZq1BlkN4JAoIsxTTqzqdz/pDGnjyq8XBxbdMtHhkHsifyVTDnn
wdm6rghWw47FIVwq3xH4CySEL6/12q0dcPAP7uG1bEj6n93C9EO6jMWdfE85z5HN
/Tvad4fjJSdvJlyty91D/nCUGzaBDirSIBX0vxr9ThoeBCYXVvgVs7goiF9bABCn
oDhmPp04JYQpC/iNhe61wbBUO9h8U8rIa6f+wYyDGy5U1xviers2pheljerm0oec
cFLLG2sfW5IZTYp66fsogU7weMmlJkblUXKwuavUzpPT4fEwkUN9C1y7UpYhHfM+
QkrKdwgFYAlviEporXVroqwZqmqwaRIFBSdX0NOaVDR29+SRkOt47lBu1Qj6sc5S
2Iex4oWi+8V4g6moxBmXVRh06ZzP3ji1Iw5mqbMC+WxtpqgT5VfWGHvjez3ifDuA
TnsvhQltiSO4qRRhjirLarnG8bN8Y/RRznFgs+gej8SPGqXNbxswRMBfkH+JzbsH
Kcs3YyV/qGXz1ShH+hg0jJ0xc+0xN0TWCiSLOefvcpAyYfNY+0Qj3vhhbgHa5G3Z
vCRnT1mKsO4nb10Uf0iQTum1UhTrJJSnhVXZegaBlSboSOT2CFpNMsUkgApipRZF
yjizARzlwY8MxhBAJgTk0GjGIZaQaOud29vix81ZWMPrU6SlTj4gEgpD64JqfJxa
ABjBHjSJ+AuvLT+rnqFN7XbP2s2qvqqphzMBx1SxXS5D2ZVtVGEiuNenfCUF0yEp
mvQxfE1ftReT6Z3Db9w6H6h4ffTZshRdozejV4RwkwpfeJR0afvCXmmHTdplPM3+
gWvz7puSFj5WJ6DFSdxD2rv+i2Shv0kdflg9B43ByuFpsQDwhrg+chR1+s41GkOq
TvpautPxP2nNrbJJxEDBq82XJHFc/SdlLj3BdPcMthtA+xb2/HeYwVrSWV3P59CE
9bkDUaAJSKdyTL8XXro3udPq5072mHryVrw3cAajkFeEeQFauFuQ9dHJaeqpGqwj
ZbJe/kJ91N1+DGBRU1ULtnnRQU/3wyuhk9BPCSIR3I5/8VpJSNc/SvZrsJrAv4MN
sVZJw8I+F3WPaA0BoKJPXx3QofrpIPvUNcIvYnbR5KrEq9ZHl5Kgtc3a1Y+Mo+/N
yYJ217moQ2qDtKKbcr+kMkHNhk8q/L8UAPYy0eDUP81jI5npKS+SAOrnBFnaNCrV
fb623PRr7TMsUKibAuVmkP9qCWihz27b2K6EkW/KXKWvlbpPcJzTEub6xK5f+GpO
4+EZktvMRE3ZXoBFgkJDR6SDJWI8oxaMzpmvmvyrjIO3YVF+SDXnnOAxhldvy/oE
UCf7PkNrnhwAlt0jGYkWD9k04FtV+FBmRxU4UpWvXjiOBaeo5TqGEp7PCssCNPy3
i2ezIYALH9JdG6JzMycx+/g4Ei6M1iHStFBbYp1dMFBPTridpQ+E1+I+kOMLSH0M
xjz33L6Sw6KEH/FpZs34qY6rAOoi2B+q7AL44ls8ru+D5Ih0C6JXB4WKZq9zUlVH
mcyjm3MFioJYFpKV03T/mLDD08bnlPbjaO/WkqvNQeBn0ugnV4JR2EQF2ZnfTQ25
JqGalL+7yMY510CFAOXVng2lPlCqV4UKd7jjeR5rWSmISVT3SfNm5E4meK+fraFD
OMhWjvmL3rP81g1scUyC7K1h/FC7u5Lv2gNmL1gPND9sS6u5V/rjiPXUuUG2BOjs
G1JEjt05GsXRU+Ux76O7T5DpvpmhvwRVsgfxdpmp5FPjMwBV5qypA+J03qerGAbn
mX6USL1czNVMbFWkZyH2lrjA7Bryikn95CaOROwK6Nhd6oAUU7+M2nJC6mdO+UAF
m3eMY7SSj2saCeBFN6Rz4IFFZyOTT6Gyaqzt8Q+LdJ8KbmIzfLKAtSN1ip0Ce5P/
9BBBQR+wEkOa15M1A5qCu+lsaleWnM/dm5T7jXush3MrCiWRfNVBIfz2vbV3/RX3
Mk/dVcqKM0wuw+KPasji7W/jvaAs5bj3kDGGmqrKv89CwXdl3x14ykN266IVlw+J
aI8Fmmr+VQr0INnXx4sKleR141c+an2Pe/k5Ng8Ydf3WtaMYwBIWdhx1ZrtHLPHO
1e5C/JJqAUERqiARSy5uxJMxPKCAFevPHv6yxTf9/dvvcFAoTgfaYyoPJhkZUR+J
73XaN0x+nMPsJCR/lmJTQuTr2Jfn5z0hJOeqfvfApLSW53oqZczuoQ+GcrJPiaMR
DhdYF8f67z+wLkpmpqwSRIRM2X6b9wF7xwL+T9znXaVgrW5xyyayUkkE+XeZNO1O
3B1GAwHmPBHIj6kI2KCUMdL9dv4Fdmq9YHi0VLIr0P8wSAgskb8UmhutWGk7Q8ao
/XafrEi8vwKeRhnAJIblDKuTtcRa9UZWJlDdo4kFikQqDF7QjL01iNwxIdxJ05kL
j+184pR6spgIPVOXsj7Qtzn4kOzAQNe1U4Wj/WG0Kv/+ynkk9nwDVXKS4KV9rr4Q
NYQqpxVcM0WqvxFP/yTaueEL4XgwhI0B4P4dv9BUdq5rUZG0BIh1KjxHIDl1kkvx
6aw2CyOSTdHGihAh7/XUET2qeOENQjYFF8p69ieuhbmWxFNCRvjoyIdMcRVRXzVL
Y7yeirSGusmrvJaKGvjzNlSMJDF158EFksOB8EYHo6az7t4CMM8VdoZ9TCyLqaPS
Uy0gItE+DMynZoUxP2Hel6jqpNtaU3LJ7fnrEKJiqk2OjnOVHHIVamGyIz755aGo
HS9XIECtxWbe1oyuQqogQfqRb3gshBvbQjN12dJfSJkJGygg3ZNKfJnVobzBaajt
615yB6xwey5fmQcMDGe25m0TI+aMFA9Hbe1bLFAlF4aeb74NCPtbUFN4+t1gAOgp
k99xGRTLt1oP21GnFPYw0/sf+fjnKfEn9R4c5xqfADjKpi7DXJPltVNfgCR1I49c
Miwc6YK0GTkujPbNZwRBRB88fvYRBvigHOEPyLI/3wyj+R7QL5VTghwbmFTigHdZ
LhXNDq5aSdRHAU+GYYlhTmngEgv6IOwKYJZBExxWk3VXKEfULlkLKtn39SkLPcua
Q0NPUEmsNzGEV0wviWvzMoe+QHIQSi/4F2S3PQEmztzqG4qY93bD5uckLJR9QP1o
P9vcwqB9qOJD32QHOF2rNyMUvbWVnP5o2c+3GpYWyiUbBFEHEH0k7zrnsm9S59tI
X2zA20j2n0vU0GgiufSeVKqXxScHigTc89Gg3h76pbEGhrnsK16RZc7JJSMjrAM7
3kgRKIs1cmtCYQ65Kj383o1ygUhot0ggoWXfIoxW2rSAnDNG+oDYo2zSS0R7gnFj
erPTZQt0tMFuPnleyLUREKmGoYzEa3m5lPopCLFI7qen34NlmDdN97QcU19lVboE
2vh9Grx3nljGDmAJll0avqLigAWbOUtml+0soTP1NBgCf0czDYz2tlf+KqDrBX6m
9UOEUiqF6BMSJlE83UqC6OGicxpSZd3cUnlLykEfmnrKUjC0XRSvOW1FM2uCEc7G
VPVnXt9FGmKffWrNkPwD9/IypGIimNRBb/6UFYZOrQd0DkRxd/FGuPV/mLjrv8xo
bm7X7Ilm7UChOQJnbTGbpfIku/elo0mG90mqzCnkgfoayXYxX3jaB5s2zUIwEfyJ
fuyrrk/vzqNME/pt2T4zTHXiX9B4AiWy8mVtNziImq6ForfhwJUGb+eqn+WYPfcv
ndPV5mZIAyNbH9duTgUvd/oZi3yl4eKpA/y559GqWFvyIR8BRPwrmwapELcaJmdF
pXiGhbDXo0KRzMTXe+vGRZmeKNl/3udHoy2Fqd4XXaBKDoHRhkwFMYThCKF+4dKK
6eX05XqdhVrnb6lRJrRtntxXQXK4rmxo6ecXKR/bO8DyVFpPNn77/BYkWxlRPgoC
e+2+rpPGEnySqELN0mKZlxIgEM8qX4NezOxiwuPtUKmXFw1a/RYmG2FobaIqGYXF
EKK/stYEOmKuA4oiZA8e2lxJ5NZTW1lP13Vg7WdZSlSe8CldyniJByIpMlLasgh8
2Eeds5BXKfBYjJe9MMROBmlmnq+1nH3+K3adcOtR8VrSBkt4LCi6ohdpwkA5RPMA
Gaq0pbsZyKMQsGjWiGr8kF9owtCr9RJqAUeT/61bZOvGK8lP7+8z0E8nzKaJyuXB
WropVVUo7fU3/WFdVKPU3xGL/EttGblNXBd4qQCcQ5+FGUCPujx4h5dqQJI1bmbI
ag72fFjzs7WeBnJ+FBk+GqXPiIVma9w2E9gr3W1QD74Bp2QITe+290e6SZVWiu63
vlB20u2MOamRpo3C6UfTknLzbSy1GlSAHkpVR11s/ccJHr7lt5rt2hQ8Ebg6lOmZ
IviL80Qpvmx5RVNhGBw+Ytwp0BMw/Ro+y4yfS2ObmNeLNzyG/RO09ZS2dpOqoycM
BA6XaFX066Jr4purzQZ8LJwOAbBgCcj27Qkq6L5hOZ6xpXywecfXqMaKs+CvLPuz
D7IKqOYZ+3JrOcnzaiCroUSZqokMgOr2Mw8IVHQHuteDBZxpSvz8ChX3Sc/Vq7Lh
GFvBcZ5zCM9jvJWvfUeeCTDmISoWYKQ1vaGxoIr33yLHOWGtfhAEVGS53liJ08sY
xndExqY/IxwXPYjS/n2MYxoF0I7kicuEf/Dkv15CopRw+I7j8k6kaIwiKgm2A4sS
nblgPADBkmBzaCwl4W99s/ina0J8LAfXa0PQ0pJAB5yzgHdwZByDZ3Z7hD0qhynZ
oFjIphmUn+L1X9YieJ3W89A0P0KGlrxiKn1qWswpfOkoTt3aGcsxlgybUb9EnKOd
KIY3+qLhaZcmbppJctN6LksVk6mzbRXly0wAqiOxRWXSKBxI+K8k9nGgpeirVs/j
64afSHSQIzhjvi4A+kQn/P0ARP1+tQgt1eDOAP4mrTfT5EW2QsPdQxvnpsU3mNVh
ad0E10U1S755zw17vsvH8j+DWxuRAZMG0BHpciCf+pyvJO+CRYF98n6IIunZAQaX
Dtc65E62sRZ/e8cMIKfNyXGcGAmj6NPkAFyNHHoLOB9MbyJJNcHRYbD7q0W1UO5o
/taiiTIjq4ZsoZcQzoYPuJotXkZ1sA8gH0ksvF1MSHksiXf//mWQB/THJIlo5lyU
IV4uRkGpIgilKTyyrjgXfQXlWiWlCiaxVXoJXECB9YLCU12G2i89PLbG4pdqfaOW
a2wj6Hzml3d03JTcW3rXdcqmhoWhZnoV4dHMsVl8bnlT4Fa7Ga5TdCexEtGcbR9a
9uKzVMixo0YOUACpyENIcf4MKrJtsPOIK0wUI8cJg1w+YL7mxtKuWQRcN1m41t2s
wjbb0fsBsWihd8JNFqupJkqpzqu9mMIGHDa3T5BzoIPBoTfywFUyyHibHhsGZHUj
pAwJrF71oh0BTrkmcWFpDEnhiGqTozth2xs9bhALNJ9kNA+ynydGBKusRv5PzFzO
n96Nk10jNPsG8kMSOVXxFfd/QQ8c+ygo+1ltxnzn/RWake3d6SUO7LHHaHmL/naW
lXX0pEyMUyofWjUDRQrfRBOogv8xEwFuywjhOe/Fyrt2NA7qEDHKmsaeVLYJmnRn
8gOD3xL6erQHS4vGiEuSPCq+1Au3llm98hzWCc4i+4/rBJzQipbGBY3ygEBbSjkd
JJYAgeWn0HxgrBtzoAKrnspu+6I6q3dnDEplvsX2RNIq6Y9Mvg5i7dr9Wp5GrT4v
6ICd/dXSFTr19+lMkCFVcvh2VbAG++vkiYmNQDUqR42rsitoRVXZs7/gAc0tmP+8
pXQJlj4Lp18qZu12q6L+kHtIzrA3mGsXE40CWcxwJV3nE8T+U7Bh3/pFwSfTgicT
A2s24KoTlD3DvDv1DVvjkcl+MWv3f2rH1bK3aRtbbQd0tQV/KsWmA6ZuUyguAav/
vKf8W0gYlu+nPzxCLfdnCND/SHX79eqaDtm7vV1QssKYEIe0RFLmStsIRVGLNZZH
cbl3tR3jLR6pJjf9gR73mgB4dWz00FOGr7q5VN+EA5UwwRUhCumw18FrsmaTst0i
Fb3VLkF018AKT4zVqjs26H3sQkNDbJ1wqgoSjT0L8RDK5U8rv5pOsjDc2VtXLjnU
yhoZUb5gP4RZ0DXWlkKTLPzEJWB0W06cMkdIeMzrmGcb7/17aaQKRM0qZQwp5qoD
Vm12r1xLPK25gQg0C2JBoLAT9/d2+EzJaIf2ll74rNPIB2s5zQeisfKlNNIHeDM4
svbH0ZqlsDunI7hqaYTwh4Phm0tBDJ1M3Qk36XdLGz1JsvZc9iJyF48SnqTu7Vxy
OribVrvi0Qk2/FVnmjKVjMgHIX/nPZd0TFh08o5bT3T6XHOqpcdNEzuNmTwmWbE5
oAu/Ba9275tUB6VQeBkfpEJYDrobSjErD7ibb1KMXAQkzgpg3cB0DZ7ntSx+0MM6
4k1d7rJG5pUMzOfEPqxtmD0FtlQDfDO978DGINHFeVMHipLPCwn6YkE+0qYN9z8O
voaRKeBkcp3J5vpP87IHpBeNyWQ6bYZ16qv3uOxJd7yN/Lx5RSNY8k7nA221ecSQ
sDOz7t18PqDskdEf0jRPt1lUPl667lL3U4DttNHg3oPK0p+iHWvbuFYxiHEWAX4G
wSIOg53VOWOLws2ym0TseSyqn9huvl1zzHMy832o5G72LsnNDCrjrmso6lW0w2c6
hg6+hH5DjIDY0s5vyHOfR/WLV5QdycpKYA/erLuNEbD5dHjiW1K/PS90IRG1qsdG
yCTm/pUwCqZwKb4SuYuRhZ6yK1RJdT7pbe+CnQdyXVo8BT0jGrwSkAHBpqck4B1T
QPwAxdIFJGUiTY70vkke2BiJwayEpHUcsCpqKBpKf2Ozd3ctD9h6yDZ3XqgNa63Z
cfkc05ln5OIsdH87roykH3EtKuNX7EdnStEbjiOO+uw0jRuu51/hhS5ws/v7YHUk
eU7XjM90pa2BEgSqILu10yLkrgnNFs+XA7MSLjR+sfFRWu4KRWuThIktJG2k/FqU
xt/MaI0hkbic7T3akoQQ8e+KnFRaODrAA0Xz0EL8D7VZ6mbJu6C9QXzwzlw33joq
PUZx+1ZtCIBFaBRQsXQfNVrovLJRkZ/XRfVQ5ZGvDc/LxrQacmlQtl12hckFk+Yn
7o4TSrN7G+tGOWEcAnlQ1z80WngKzTvT+UXK6s5tAB0SPCs7earJlMXNYBY+tcy6
uWzz8XPqTXoSIC5Ql8Fj5ujOU0SEcBSlnnnLByaV45OXKTxoxscClqKEsl/546P8
0bvKNs6mHkQG2ERF1kLgrriclkonHKLvFJkzCvn7N8RhYQ9hxqEZto7WvG/Af42O
zucYXaEDr/Is2BY5LmxAc9nUE3Mg3druzWGj+j6mJtQ5A6R0Tnr+a/fyNFONFL43
6hBXPq3Iaxp62MWkIJS8DYHR4lElkvQyPgx7XPwER8zNZQdi2Q5fR0TN/jOjpyZ7
3a/ZQewqW7+yv6nDK1dDY1WkBmYecf7tNiuBvorVJyrrjwGXMoh8c4uVcniS+43V
B2KbIfAldwxc3g79x7SrakT7MhJSPOoZIPHpb9kqQxpDMOU1RZ7l6i+Er9NjjUi/
WEZY/onTW8SUKUN0AAFqVBXGWLb0cl+eRTPR8lVTa0idL71uZmXsy3eDq/imslYE
nA11+cdixmxL85n4QdaBzscoJHOv1E6UOAbLu2+wgUGI+XPJUHC+QanN8TOpDL5L
JCy6+DJoN1jImQifCYklD+t29Fu8NfUGvFlviMmeST9sxeb32m/kM3g3epGQa0Dp
rRapssOgsm912BeISDpHrdwl1d5Py6vZbnUN5JOVVrvPNr3678xFpr1IGJAGnhhv
N0Q0Oc0XIPH7F9GJkJPFqk5wU8hsSgq29BRF9UBVArnmmo+WQGfMDi+t7Wc4Idim
HzP9YJ/X65kjjczWaLY8s3DPPR5yoAAGcFNKA19+1bi2p3Vz32BWGmvc7wvqHHXY
p/ERZDWnnJXsWte831Sr4999jmcepO+Dj8YBcSVS2aOd2dNyPQQNTnyf4XGh/RZK
goSzxKFfhi1Ju5L01RvFphNU10L5nL7LPZSOaC0vn3J31D3Y37ezT7wUJ05p3kVA
QNPIN2CtxpQR3KKAmvQuQ7Q/INm1A7m/e+1Shuu8nmmJEgwac5dyyD8cYvVvRzLp
kFyL8bZlMcY6//yppk4POFA49rjdGyfFFxdb+hVnDJonWIJaa8NsWnvdLeE5kkXD
2ZFk2XyoUMOd4jvaEuQ59gCYuLNQI+DVOeYp6dnoXcy1g+308x4ejJ0Vy84P9LgB
wdeWjKTgRy47dL2U7/syQueuMXNXNDfRRe1IDyoEBBAx6OwT2yyzpY0ehhinufhF
JufdLa7fUGOvx8Wv0dHA1I9m21WCABy3ZYzW027AniqTktfj8tmb+FuEsgadC2dS
at6uA/1LL7NFcQy+YFynNOI57HNkDxWYRhGxboCmyoJGB0wGXBjH9MxOmNqh/Qh/
mXSMBbcXGTe7V+UQEegFzd4k8F8jpEFJ8728Oo+JNiv68AzVdn40jlAvVWsw9E7V
dNt6VvWcxlzvCvmpnMKdZTnRPDJX9xPgmqUK4Z9S+QaQbQD4VrVLtwyh69caokK+
poetXQOy2q4Qv311gssWBM4f5fxDf3ShEHpw+62xPqVAy2Z27/RC/pncXkUqQEhI
8EO1zcn+Y7nYJfVKvXsI05b+rdgf37M1LCmve3Sl0CWkyPg8A6O5R2OyWwIZRLIm
l3K6ClgfkLSutHg+ijVTRz3ldL6BRyWB174il1w1fE1r6bseiRCjY08WYojiqWSg
ap9BsNsLshmEJCFmkvArlPC+henX/MxIwM+LC1zoTyQAVw4dvUPIrbb4b5oCKMNj
4LT57u5f8rTdTgiwhH5s9JuIkv98DPRH+al/u/npVp143MQw+JRxVWfx5H8f1dyu
743YD9j130kdd+/gpXSGzbiR1KqFl+aMCUZcoOg1T9Ug7eZvdcAvTeXx7GVPtCaW
q9UstqOq1LwocV3Ryx8+cfPvT8CmR3nOpTfT0wC3k0bT+0KS9KdzLwty6qHPjQ5X
cdjNRqYMTO/Juw0hp0FGHPHfHVd4WonnRhy7Vt0W6bdLWXgtmSReYlnZ6zxqLRer
YFojt7Z260hh3w2z7kv/h8r3vx43ohxIeP4KgBvTSvihDSp14mvoC22OUvR95AmX
3Zx2vzwnzBpmexd/9zeqmFOtBvhwZj+T78ho+BBFGLjR0Ph1PhTk0iylQlASX0vy
mEFrd0J9st2idFNAv6RheHbHMXWRqdO2XwfYRytR9oopdFVW9kcP8+5pglAEg90J
j/ft373xMjoxMHhJ31V6tBbVEdOzW/CA7uWqRoB6v1qy8h3kiOe2jCcwzj7MnYq4
vS/WqVM1d78Fmi4Rs+LOZuApnxdA72YTcBjjURPy4lVxLZ3//Guo1H26ukskb4B6
xuFHJID4iMsI7WJMpD0O8RVSGrhMyWmuvmkx+BxmE6goxqM6ZPztJkzHWqTm3+GX
86Qur3a0jTWq5kcmkVFqirsAmKcomOkEorKkRHLKHRp0Gc4K/EWT1u6EzODv2Xyl
LJoP06gZTXKz9Ce71UIYQyQRjAVu4DobvTyaKY21ilTmMVGe7SOq/hYGDc8bg/cA
daLa02mlxdZb/6iodQH8Of92DqdUYEzJlE28xEpWiZAC3BEDtwkO0O/exYgfjEjS
zAo13mFT2evQlKPkFEBCWp0dn6NnAHd8AuO6WgMbHyvU5Jj/VmWScr+onXFZmCcA
Wla4KAtZNIEuYbyNXJLKZvlQIP14bZ4emeHN8O8zNDibbkvqIORxRsohS1op0V0q
V09zGltErPbfrqa8LQZi3JnfjM6atoz/hNap9I5CoUeml69dX1kZbJfp4nkOhJvr
0IKF/TDu+2Ju6ryIdvHHhLw4jZocngyxqHc2mY2rR0I8bTH6CMMQFWsJpEKxpKNy
SL14qgVljqmxlf4TawxNzm8oq6Ay/sr7ASAlSWqqBT7Xc3hVSBjZEBuPzsYnfHsb
DLh45VE4DSQlrLMAQkB0LrbuoOFDy26JcnIjRY1I0UN0ZKDb/8SPAgk4YZCf3SRN
ZfxBH5vm+3Lmum3vwFXL+d8WVhb5nZaGUFpUi5wUjCRqCYOBHwgKAq99yoBtFA7J
5qBbE/DUxr4oz4lRljbe6OA44amjpyrro5/lG8tcMXN95irwWzfmtdAwWG7vTDtN
OBr5NWjFDD8TJrEX1RBAFSlq7YbVNkXxqTHrtyxCPHw8LxZINoc5XM6nJy/t8jDf
KkVwmLeQ/FGmNDeolAlRl4PnILiLNCxqdUloh5xg1QkG/kJt8RWlyIa2lJfX3w/a
uPVp1TjuZ8WmgRHYZr5/aXbkIiY/m8/b6PGzc05lJhg3ohU4/InMYx3pK756uoM9
H8YAbwwSMfx+qsfnP9ZkRulRkQqYNoDxPU24svQdtysYgUx8Sv2oBPv5GXJh/Mep
6mUMvXK/kb+hGRCfTcwhyLcWgD8ap0h4x8RwftQdhQ4hBIZ5XeAuPftOwWn06MxA
J2tOFsA2c6kzxUYQqiZ7bSgbCEl7FwD/HrNpJxg8zzCZKCPuI1jBQkfIggRfb4+1
01RqnF/+M9D5y0mDsw4yZq+Eexbi2x45WbITJqO318RwO9wJ9YXGTCadytTTo4hl
3HH5IJfiHzhozgQAz4O2BEs7g28UPbWZh2bd/gRUuNwHBGLDj3ssak/+UU5HgXo/
m7FmziEiD3dYDkAEjJSjnk7MZzchfvsFpdnAIy9J6mpxujF+svoi8IZcV1G/AX/b
zVuJx6XkjvPTGXgdk2rBWoj1E7S+6aRjJLiUheHzX610fM3k13wJouTijMgYFF/S
RexiPRYHTzYpqpvwgADbbmbRr7/m7WUdrYdXOKAPR1V9coqCCcety7Hj232j3svp
XkWyTQO4BViBOKObJfTrWJmzJIWQiVjj0KCnjln4iN/EFd21bVmw/7SrGQ/SRlwh
F8jP2Ji/M0o4KdsxrtjLVrw95bSAZ4GeU+0yT186wSZNtMMLnf9HQp8NvkZRU9Zi
TrE7Fw2vWzaxNzETcaHEBfDJYeYiNv2y56F7JWdArj/TWqLNBvtSIYcG65ezIlex
fzgqRpuB7zs2lTHB9nImpKAgSBPUEVh0MfOWrPIJyDSWoERms4TTzkiqEUTRvkia
n0PMaeZa+OZ/mlPqdpKtqKEhCwkTocM2kGrqO+NIv9mUcW117SBHYsAnUpjmHmGP
Mz6G1Y7fcoU66Oui4owA7ZZKZpf1uq/d9WZmlKu2kFfaDlYJXtRfMIA/GptteWLy
mb+gULUF4my/VdHPYmFlyn+2+tY/tGS14EUg9PNcndcJ/JMKv3QRiOl1jjGSsU23
CsE1rxpNSNlCPY1gJo1jki4BSL+sJVOWQSVW1ML53DHcdj83gpX8Sgyf0xS0upWz
SFwla6AhZXohPKHyr1KgO4pVp/vMUH/FJJ+Y+3Vh3Crxr32ycn6uqdPWnoJHBqY6
6r3mnjPMF6Jqs5Z6F30g4J8G1cpeMrYTdsKxk+XUCze2JWcUL4OnI7Qh7nE2T1fI
oL7PkiiBkk4Q2dz0N/kBgs+6uioGWqd2T1qZtPvnpSNu81kMtAXdQCdAnq20RN2x
yFWg6W0YQtVITc+tD1kKOYFV+U1gSseHOsHRbRNdy1BLUsOTPHCfi1LCYhGslZPf
9egGAAjDYs35scmf3q0SKmFU2u6MGc/6PRgKcaM4eZP4Kv5kHGjH1t/R3enIkmCp
`pragma protect end_protected
