// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:13 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LeYx3Gn3KF5Q1QMveNzr86Z2js/aP+39ztIaF3eCT2GPMYnYsJXksBJeWiCpVsv6
rWNSe/go2LhPQTEU+c+OciL0HK3P5PvpV6rXJTNozCPcRMG8sh8TawD5kdGSNU7S
YOlwxOSJfWMUPjN2gegPLgEt4YtuFkc3O93ICfx/atY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
VluPEzJ7guXpdcxCc5W4LddJgGXflWzMyqG7XbwK0QwdPw9yYtbn3+KJ3QI84yj7
OqOZUxPA8kLs8sQtzXFyB4jOv4ZzJDnqWS6Sm6yi+OdbKeBjGRmG8cpz0tN6ooqj
TKzA/t0BF6vn4XrzSWw1Elfw7OFaNDn8td1xe6r28pwX8TpV5rAcWD1MbZPNAyRV
ngbGoadfod4/1aEm+Bazw5yuH2+zXK8XsVyuv7dz3xjeiRy7MwXjuafS5dEAIPRf
fenwh4N+QxZqW0MxW0A3V7cgACaUGkDG7+jHaGMG3ERDQr3PD/67IWE0TTKAEb8J
6eBT06/BR2JE3zm+fctDJf+jOlAKxG4DT49RjH5FEuybQZK6PAEdU+JWWh7BGAN3
+BFN17ICl7x/Iny5x3MoYK5H8cR7Ux0X8Qftzni7ZRdbVYP3QAVd/w7fDXmYFnEn
OPnwloJd3IK7yDngrZAQyJXKoyuF3DD+7WanOxsuVn7zy5pDIK7UT4bpjokoomXJ
M7YEcbs1lXGtqdokcqS1zYe7bEvbr+34/hvbX7/b3HkUcfwhbWt9AZn0zNF/Kt+B
WQxPXSk9wd6edtytBmTq6gmWesDPEX9lC0PSYyVVTsgg5gcEycKGRE48ou3sq59h
a980Ic0C/qHfYnVTMYu9gzu1+24t0IqkDnhLmYSuB7brEr/gHzEB8l1pnXjZVBXU
2rwQ3Eq76UGNOWbdSByuFpNmY3NaCH09Bkh5AhOaoos/ZAd4CESZLOSG2t8WPrBp
0xDS9AVsj47o4R7jTT+hCKlZ9wdrL6GgR//ROZ98QGl0WFUm4rl2byJfPXdhfYr4
JfgKqhwiSqbsUACF41I62dtY6W6vHfAlOS1aL7gHBAHJ0x6EpDMQs8XDeHfG4tP3
mvxOScGJpEY4RiBUwAsMSeQ+j2/Rk8w+7pn2jJBGu6Ez4sCczEz3+tGSxajyy0Mr
FanPUFJzLLiq76XMhibZ3XWiylBmi9/VXhB5DbZ9RCkgCCdU1vKrBMPKNT/M31AX
SVesZGDu56m5etotVc+ItqgzS69SehylG4Pc8KgLhw6/N0FPIDI+QkAlYFxnof6A
Plyv3Vw81QE8N2s2Rh2YosSsf2rHkA+oF2c1hHRzehTY4chZRgEBPHIUy0RJjk6h
Z46cu3vTee5LXVL71kb0F+dyLxb6BHDrR+3KrU9+0FLJyS7lcFOQRqWJboXoC429
q0/5Vvjm9TDpjNvas85rACQwDhlvbG44s0XaqIdPzgukIyvF8Je8rkOBVn2xnyhO
N4Y3MN7+kHaTgKlQOKS0fmRKAZ2vnfVnbukg+mcHhk+6OVy/bGstdxgFIzZzKbEx
IDpq4wDQKI/OnHMQqpHlrLpCHbZyl3drWa6gIbxr74nEqx5Q5pcwU3awT362wr3j
SAW69z9L/1PlOs4MuzLXWLwy/iDGg6ZhvgIO9oB1iVg4Mgb/xhTv281VT5ShuKtx
PtOW8toBXQk5ny7N2jhWGKCMQKJwyv3xZnLxCefVB90itUyk3/xLA+nEnAAuSyph
jaRxnC8sE+SaCmeUxhfbfhLjg4d4xsvmVI0afXCk450BoMpGoYJixhxBsRreThI6
JNo8+dQFm47htx3UXaoUGgHsEa6PGZSCFLnM74D0OTkrk0bjkZ/Y1RRTUNOYYvaG
B6PVv3y/UwaxnpJDuYrSlSx4wcLN4jC4BnocRI0W7ZDeMK19rvxJN6yb9tNvkAhy
ygaFA02AAEcbW++LYLyiZA4VbNncIB2Pp5L6/7cI/r+vKTcGccWnmHkx7y8OvW/D
OIeCPLzgFSW5k8C66soJxefRYdZSIojABkxy4SiyFWG5copuUdatZL6Hl/HBI/Hi
0xUHS80rAdREALzJ9OwcKOFkWD1KMggOZo9fZssF6l+2d2JDewSAG61brDQF3xIW
5eNYuULeiXPU+rcl2aP94hgavhEV3yK4RlKR9cTQvfMzXUK2MMGmgR8j1hcth7ZB
YUSVOcnh4HpbIKo0aNt3gaLpN33lKeBk7wIZRzfE/jR99gEeobi5cr0g0dm+lESf
sl0u1sPNQRq1kUIPFuYwv11ylZh6Eh7smapprEmmhbse3ygegfjjZ3m28b1srs3z
GIs4ymOCSVFWnIE1MjTxTsWLCoC/QrNyEkLIjlKalp32471LXZyRvIWBWJXM3YFp
4cg1OMpWR0jSDYPtldtv68tWZ6Ff1/lHkAjpd4TODSLt2ka7zbExIjysK9iH5LVb
k9kHjMtvytz+jCPEf+yPEr28uKBJ5+eUU8KCGJQQGEZ0WFQKzcni/cwDw/qRWMF1
PIwexh2OLJqX+2AvTnr2gplBgKQDFZZ735hAjtVBpcB/25qhbkW6ORPg4x65mhcQ
qzrwP7ilh8r3yGmUnZaTlMWRQrN26F6c+7HUzAuI5dYX71J+N4+/7/9StAwjD/SI
ftQN/hW+DEU0DBuChhX+QkTGwid/uJuNIdjQIGMflSgd0ZmvTGKRtsU3gaRytkeH
gYA065fjyK0os9xfF0NKHljGcls6Z3MsBfMqx9EhNHF07w/Bipk40tvobpKAecpt
H8r0S+AWNcFFv30o/ve4M6oo22hOwkxqsnRwJngFX1scNcNBLrdjstbD+NiEnA3i
AEk2MIUvBW0lZFOXrtVioDBoJAA6gINWiCmxpVDbUCqpzicfbqQF3YGd/MSn1ngT
7F04leoeX7SsBQLO0branz4lVaEA1M03kfVcwf4wU6wbKMV3bJmSdfbBV68nalwv
0nq9UGh7uZag/C9qRrzSVmcB3s2Ui2HgHBI41kM7APQ4ljL+XAq0ITYjscS5h+VJ
V9r+AVap7/WAJ5MdF9SLfCFlMWS00qHulZGTCxF1B8FcWiyUYkwaettvfzlo8PnM
nacLBI/0reL+QBHSDuJ/9GnomUPNMejfiA3Ex+9nGnzbZ8CzeYLRXtHl8N9Gaj0B
85jzgbKh3AJS42LQtNMEEglicXeGKHhXLg4wc9unZSOgYhSkeH+9QBYuErG0W+Om
RIQB2sEICVdSEZxpxigpL9ja+9C9bmPdZvPGoO5eH2EhLcSLKGM7PO8ClboAx527
Ma4wE+L7beujyqXKbOQcax9DKSDDzkS4xA7wKMEGuhoWMPfPOQLY5PvpWBTvEte6
Xq1wiXnV3o3uPbsmLqcEvGiM9Uma/dZ0RMIcJ5RTf6D4I2itgh0S0LqnVsmpcDLR
/tdYd7XxlQ9R5n8OBhgGfeMdkDJQq39NxCvlInzpsGAtU4MgRTRxgoVWLsIu5R7E
E6Lvq7qdHOzU3zIpzr8IhfTaZsnIwfSXnwJfh8/yCLSe0a5A/AcXZuhKsnj6Yidi
KMXa0+Mi62nmcWUZ9Vv+eCuWCE12DeemNWwYZK25H1Usjo7In1sUnKvY6HTXNbUj
TGJU8UCE5D32cIKrj8+UQesaDernpj0PcJrEHBekl+JwNSow+LtPHy904dpotKAX
R/kfq/Yt0y6wsgKYW/LLcssd/07U/l5DuxeZdIvpjlPIXDJV/60rf7vYBgqBRMA3
xX9363OAJtG7e7Ps4h3klk00kq5zRibp8dfygSIcVpdo47Fx1vDJ9wcpvwswxV38
j02jLA82jEMu4W6K5dGynT6DeADBwVuq/3Qex5gv4Mz4K4Bth4pY4h+icjNRuqOB
sZtUAlkJuDqsaM1IdVaHDwBiHrg5dq+qovpCqXFpxb/NCbWl5I07G0yXO7T633fp
CK1G1NT5o/KRExsVRXw9CR8WltX13wE+d8aVrcgAfj7aFBmpYwOUJrRFgERdnXDW
vjjbVeh7/EohwhNKdfwsZV5pl4pqzRnhYP/Fd/NWXoJm9gqjHy2ObRJHa4k75H2L
l9qyPiRE/aEhNIZnD8Fs04YC988Z5eepE7foHf5ubaAtaOJgDUg7K70uCY5m1GSA
weeLY/AbGjhVSj6nO3sRCU8K1lQ+CBx+Uym5VoJ6JBuYa9c5d+3O6WFeGw6HwOQZ
7vXMVGPrzO2iZNO/kxvHLT2LAiuZwr6M9tn15EYu5yNhZow2HglWwsRT0oIrEaQr
gLVX2m4+U42BIImnicuNNsf/Dw5HFCVZouq6yGXWFigSUWCDhnHsfmk2xbNxF5Ek
ghwHdnUcwJ3K68uGyAsLKd2vtxMszx3vxvftgeRDdX95VkfMIN6Fk99xFcYreJO1
VFubvdfF5ozBNVu7V5rJfbJebDTT2XRTtYAKSLzEOIIDiAqVu0Hku270DF4DCQBU
/Nh6qdWhlxIJ6Kj8hdI/FBoE9tWw7FdeK0cfJlBe0o1hRTXKvQZHkI2FgyrIdqXs
1t2M94RsJWdf2sITCMQbx5lguvURIs5oOrRwBoNVWAedv/GdERCV9LKyTVFIFydW
Jb3u0sM6W7kPfQ2xGf/VFiFdEOLv3L9kTFqk4ewSm+kJwQZ4cx5urDznHYz6eQ2D
r18IFMfzO5jgG1oiep54JKwbAWXRBmDIpPv2Utu2rfktNvvaknCSXstb51e+eQSJ
X+O45sPwsHP8h9APekbmsLJEcOHzpQP8guWt3N29wtjJdkQWcD7p/2egpvlEqPik
LjqOL2ZNtoT63GzaQWG1TAuGU/IjOEXgPsehlPDkDJ2RnuqtF8knqDubyRMoSkV9
ZcG/FduH40bpRA8adsJOZL5KaujP8xtmEfBuvu1XjUnijoQod9AawnMjWKJTrudi
q1klt1r9gn0/cGob2/HqdoLjYRASk54Parto9JBDCrZ2eZHammdq8AVQl4NLe8Xi
Qif0ZcmWYUpP8ACNQwj5IOsVR8lAmZTa7BNAERttr5TKqhU9vfqL7AQCZXth+Jav
ZqE6kPtrkaea7pUArcyBAJTI9b+0uc5e1u0SfJ9eaq1vpphr/IBRw9/nH7j+n918
JUaIpsU/AiwyP7rAxmDqpDHqOFOVu29tEF2LTcX4nY4fvn+xUYLQIXSyjVRFB3nG
NMtyOrZQfq102rPO2J+XrjYcektTLWGoTbHosh/CH0l1053E5ZDx/dVEZbMrmfsb
m2U41Qdwt/jsesfLKHCs8bvnuV8OBpXSp44/iNuNwryziUZz8kOaaqBp+ji0XlJr
ybG/8i2hv3rEz5c67MyMZDlLmPnFQqhYEDJoDjKtPU7b4fejXIm8ffSkYwGz0mkp
cNFJkXOkV+SLis/zjAhZtc6iDGuiTRKsFVcP//q+wfL0OC+e3vx6PuUoaw67kyFX
DeZUbwopP5Gi5nYd0ud0F21WwaNCcwwSSIsILUm2k5Dj7XcKyiGFZsCMHAkv/VK6
2Pw4n+lMe9AgZ9DFAw7bjIxgy289egdIjhpwAfeLACmF/YPjoqSTUv2HIxLDDfoD
2Q5RpcixZbYvfT8Kr82+yyIFZdA1ZQhYx1WIRhaSXazP5m9rgFIN6bIDZlzDCLo2
ZlC0CGuKoSbbHrD6DBW6D+17MJlv7GJiqZwADZzN9BKdY9CwkRupbaPd/i0hjt0u
UthjaZgQfSiISy2Zo+TNoJ4UrEHvvAv371g3cZravExL8ka75i3pahGZx4GaWI7L
trRvsx0ycHJM110LjOYxUm6ETb91zEoVlk5QIPyWLRmczLDF4jqyv2Lx+2XbtdMo
q3tY+n3HMNLMnSP2IZwU9LGmJmbaGYpesKhnRNV5MIHCe9k4RpRYhQqtkhgg+XRZ
kW1GPMA0fdvsmCJtNeT9Rz42SrXLt2Ve0/jr3z62X9wpc/QG5P6TQNf54WEEaPJS
srSZ+dqclw7wSzZNyjVJmwBY5O/U5cYOMwZdMflBkll8aejFoxMyiMwr6ZZ31Cca
onLIn4mTqbxCiT4HR8Lf0Dq/XO794R4nJDmSvGWhDb9LSgpFFmqCV83eX1knuXS7
z4EglQ9JrmOkxxEq9dc5ndVCZUGRKzFUqrvZZZEKF/p4eGfTfVvMaXdq92Mx26RS
QjdWGb29IiOSQbst43rftHghJr6BwhK4E0MEW+2slg3B9Qbg1Pk2dwcu8C0CgPL8
wjJYhB0g/tKV9h23gl1DsZq++Z4MQsAZRF3l/KVz15husKUF3rzoqq7CXVoiq7ay
dtGIsU61XM79VQXn26u1054P+gsMQj8dp9fIpA0MyYOzWGhsncawb8lU+C8M7HTe
HUY8ShORpcVquEyMo4eg+hck+V3PtQn/UPzrzglrHQkB34UpF+1hrqyWmWdgZN+n
UYobT3CWHYwRYVBbCP839rzio4eyiOkPTlmQpNhva2hiKPDflfdBlbxtcnr1o5B3
VSz/YRd0QWIxtkF6gkBob50KB9ZQMDtHgiVuVZhHTewGM0Hc2Uac69da+xTxf9nY
Jkbc1IHThgHi/ZT43ppMgJZ6PTtZ8CrB8656Df0y5v99Xc7hR/GnW74wZErBYkPZ
o7R1sEnjaKdpNdflCC4FCDHPVgcVly+zXUDP2QQJu3bBVGQLo6mn/wBsVA5hpp/d
gusYt89oU/zsMPbUv3TIXkvUJYzVKjMwHDjpYzXzy/4l2tS2xpOMyUzI+nXdadJ1
S38b6HEwcOGGbdSp7V/XlUqXnYvCcAWREb9E9lt9g6XezejM5GXHf1tyczbdgy05
R+5RVYPrAP5DsVwP/CLj1p+SNL6hDaCiZfLP6a5dEg7e42eI+6/5OzueNbbFiNJO
Iz7oOLA1rqEvmrNnQcTxfDAy+qPXPfhXMk+gzlN3a14U2dToRkH2gK2YD8lskuCg
MEBbZvdk3XS5FnNvCTMK9EV9EJywb8ZpnSqlYLkPubvBdirr8aYRbxo/zs0lIL8b
xnGpNeFBhOYTUCoA7VdjhVZMJeIrSL2JmwQ5qpUHjY+/EsiyzzJBXFjf3uQkSgdJ
utVs7YxiAohwZwQkuOGfRQcAaOENB7UVIAcDUfvj95uO0cKLDkENreXGL3hbNm+M
WRR1EMHLPzGl1BBF1DX2t+hYceSwj/PZt4vu/yOn6XUyPJaG2WyPFWppA/6dQP0u
oEfZMReyb8WQUVZTDAOq6/ncSTJ7/E6AraadgCEW3LNPPuwcAA8wzTQya5egyPv/
QXVEl9CsfX8g9DSXpz0Sedc7W5nY/LmtwYKKMVxo8qIkZifNxuRI2Yb92n0BJdFm
Z/kp/YlgmVxTUmUFOgyn7mJyGGfgyMz36KsXSr8mw5/KCHvWMtsVIsB8NJIQyX3j
ktY/kzT2EN85J63+9CGLzjAiH1mh1BkxGeXrSa3TwLVDs0vo6ADnPxgbdoL+IdTz
2O2pWl4asam2zlC7hZE7B34v1arcUaUsOWSDEbeH4uF4R+7iiXU4TpfnCTT1ieLV
940raA2hQ/PrXd4ElhSq4Rp1LoU2bOb9oirqx8456GhiGKsrR9jvw8pNoP2d6lrE
N+eljIC6e17WAa+zBS9wp32v1KNppilhq8IqGMtN3fqHoFpAdOQmq1UuUQGmrYHU
7wx+V+GG/BR10/R2nJ+KRYRSMiBzYjzj1P4AYAZBq8x/9JmaX/27wGFyCn+3pt/K
nPs52yMyuqiGx2hczGkQ6MT8eKywb8qlYuGmLx/R6cSVyPHgyEeOTAiLcHB6qdwF
jjb54Z3p0zdO5OfObS69BZdQrOfIyIfAO6srDSPgWEXPuIxnz/vTBTpbYJ10L8Kh
RNgkdMOjt3JqWbG7ZS3zCQbv1f871MfJczWqVAXinNAG6iYRXD116YyurhNY2oIz
k+oGNCsUPoC0/7kV0YZnTmPgmjU2CPSMA71TznPlyERR+LGjBOFVQ9K2tW//QLXH
DKNN8XBsFtcGDciUsdJYAu37g12yu1e4YySDTFca014=
`pragma protect end_protected
