-- sdi_ip_ii_tx.vhd

-- Generated using ACDS version 15.0 145

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sdi_ip_ii_tx is
	port (
		tx_rst             : in  std_logic                      := '0';             --             tx_rst.reset
		tx_enable_crc      : in  std_logic                      := '0';             --      tx_enable_crc.export
		tx_enable_ln       : in  std_logic                      := '0';             --       tx_enable_ln.export
		tx_ln              : in  std_logic_vector(10 downto 0)  := (others => '0'); --              tx_ln.export
		tx_datain          : in  std_logic_vector(19 downto 0)  := (others => '0'); --          tx_datain.export
		tx_datain_valid    : in  std_logic                      := '0';             --    tx_datain_valid.export
		tx_trs             : in  std_logic                      := '0';             --             tx_trs.export
		tx_dataout_valid   : out std_logic;                                         --   tx_dataout_valid.export
		tx_pclk            : in  std_logic                      := '0';             --            tx_pclk.clk
		tx_coreclk         : in  std_logic                      := '0';             --         tx_coreclk.clk
		xcvr_refclk        : in  std_logic                      := '0';             --        xcvr_refclk.clk
		sdi_tx             : out std_logic;                                         --             sdi_tx.export
		tx_pll_locked      : out std_logic;                                         --      tx_pll_locked.export
		tx_clkout          : out std_logic;                                         --          tx_clkout.clk
		reconfig_to_xcvr   : in  std_logic_vector(139 downto 0) := (others => '0'); --   reconfig_to_xcvr.reconfig_to_xcvr
		reconfig_from_xcvr : out std_logic_vector(91 downto 0)                      -- reconfig_from_xcvr.reconfig_from_xcvr
	);
end entity sdi_ip_ii_tx;

architecture rtl of sdi_ip_ii_tx is
	component sdi_ii_0001 is
		generic (
			FAMILY               : string  := "STRATIX V";
			VIDEO_STANDARD       : string  := "hd";
			SD_BIT_WIDTH         : integer := 10;
			DIRECTION            : string  := "du";
			TRANSCEIVER_PROTOCOL : string  := "xcvr_proto";
			HD_FREQ              : string  := "148.5";
			XCVR_TX_PLL_SEL      : integer := 0;
			RX_INC_ERR_TOLERANCE : integer := 0;
			RX_CRC_ERROR_OUTPUT  : integer := 0;
			RX_EN_VPID_EXTRACT   : integer := 0;
			RX_EN_A2B_CONV       : integer := 0;
			RX_EN_B2A_CONV       : integer := 0;
			TX_EN_VPID_INSERT    : integer := 0;
			IS_RTL_SIM           : integer := 0
		);
		port (
			tx_rst             : in  std_logic                      := 'X';             -- reset
			tx_enable_crc      : in  std_logic                      := 'X';             -- export
			tx_enable_ln       : in  std_logic                      := 'X';             -- export
			tx_ln              : in  std_logic_vector(10 downto 0)  := (others => 'X'); -- export
			tx_datain          : in  std_logic_vector(19 downto 0)  := (others => 'X'); -- export
			tx_datain_valid    : in  std_logic                      := 'X';             -- export
			tx_trs             : in  std_logic                      := 'X';             -- export
			tx_dataout_valid   : out std_logic;                                         -- export
			tx_pclk            : in  std_logic                      := 'X';             -- clk
			tx_coreclk         : in  std_logic                      := 'X';             -- clk
			xcvr_refclk        : in  std_logic                      := 'X';             -- clk
			sdi_tx             : out std_logic;                                         -- export
			tx_pll_locked      : out std_logic;                                         -- export
			tx_clkout          : out std_logic;                                         -- clk
			reconfig_to_xcvr   : in  std_logic_vector(139 downto 0) := (others => 'X'); -- reconfig_to_xcvr
			reconfig_from_xcvr : out std_logic_vector(91 downto 0)                      -- reconfig_from_xcvr
		);
	end component sdi_ii_0001;

begin

	sdi_ip_ii_tx_inst : component sdi_ii_0001
		generic map (
			FAMILY               => "Cyclone V",
			VIDEO_STANDARD       => "hd",
			SD_BIT_WIDTH         => 10,
			DIRECTION            => "tx",
			TRANSCEIVER_PROTOCOL => "xcvr_proto",
			HD_FREQ              => "148.5",
			XCVR_TX_PLL_SEL      => 0,
			RX_INC_ERR_TOLERANCE => 0,
			RX_CRC_ERROR_OUTPUT  => 0,
			RX_EN_VPID_EXTRACT   => 0,
			RX_EN_A2B_CONV       => 0,
			RX_EN_B2A_CONV       => 0,
			TX_EN_VPID_INSERT    => 0,
			IS_RTL_SIM           => 0
		)
		port map (
			tx_rst             => tx_rst,             --             tx_rst.reset
			tx_enable_crc      => tx_enable_crc,      --      tx_enable_crc.export
			tx_enable_ln       => tx_enable_ln,       --       tx_enable_ln.export
			tx_ln              => tx_ln,              --              tx_ln.export
			tx_datain          => tx_datain,          --          tx_datain.export
			tx_datain_valid    => tx_datain_valid,    --    tx_datain_valid.export
			tx_trs             => tx_trs,             --             tx_trs.export
			tx_dataout_valid   => tx_dataout_valid,   --   tx_dataout_valid.export
			tx_pclk            => tx_pclk,            --            tx_pclk.clk
			tx_coreclk         => tx_coreclk,         --         tx_coreclk.clk
			xcvr_refclk        => xcvr_refclk,        --        xcvr_refclk.clk
			sdi_tx             => sdi_tx,             --             sdi_tx.export
			tx_pll_locked      => tx_pll_locked,      --      tx_pll_locked.export
			tx_clkout          => tx_clkout,          --          tx_clkout.clk
			reconfig_to_xcvr   => reconfig_to_xcvr,   --   reconfig_to_xcvr.reconfig_to_xcvr
			reconfig_from_xcvr => reconfig_from_xcvr  -- reconfig_from_xcvr.reconfig_from_xcvr
		);

end architecture rtl; -- of sdi_ip_ii_tx
