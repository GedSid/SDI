// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:36 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
D3BQjfgLQt0qSQMrElBEKgjEfS8RcTiy3IJH/qFEbcXDyYMUs6+pdb5MP3g3aYBx
Xs1/w1MJZNYDQxHhcQ7fMN/hNlzwfGF7XhWYh7QbO82Xcmt6Z0MUABElni/tuG0L
/PrAsuR5DtzNIkm3GqmdPsEGvsulilUM9ouoBNS1Dws=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12352)
qd2FnLSJqqn+gmBae/d18neu2ox5gj/GEVTsqJ/4vaePzNSilWneG1+oNTGErLyP
JSMAwiWAqa0oBaxfHXU3MnQq2BvyHXZ8MnReGg05cLlvkHYO8eycJttNlTP+nrH2
Ko4gCsexChVs2U06gLURoyxTn3uSuXFtnvBJzoljC9TPuCbEQZZHSPNo7/EDisl2
+JBECmKcBKtaEhnTV1OgtNmnXwk+Hn267tMufi9bgPmtw6U+hDrM74t/YmRG+nWC
Jf9VOuH3Ki7zFSDkwWHm9OZBU2+CZfi18f3urTYESC21hh45Q3ihc9DrdAHrCybM
NhOQ6UNISwrDolS1FSHSitUQ+cZ1fXbzvkRe04HljUGem5EiNB6Hf5VxlXrcq/Rw
wOO9M1A8ym+iMbVIT9gFlnCKEdpNVMYkaYqi9kPWofR46/JEKIQWVMPMlxz8/YKB
4mVt91U90Zx5wW9lWZXoPcnZaKs9YxCmnN6hwtoFgxwY0OXPzigV/kTiMlD4q0WT
uC9IDWqRXP9lrv4SKFX0viGWI1nWloWNTUeiCf+Xw/f26+soiAo6gMQocS25XwRr
JDEnMyLWAArPcnH+jbKDk0W6lvFNE/REDJ5nKhWtuGNLFgy/t/ePdrgbaypx/wn+
lc/L4h1A2Lkf0hMkOWsFuaJh1MVz7byQbVL1HHOaBoeGY9yYg0Zm1LbbxycWvMpE
dwttt1IXLZXxZ2H2WbTIdhzlwibLltdPtAzhIu5b3O/8nq2ZU4Iv+4ZCLDKe7l0E
8i+79FPvvUMdxMi4fr6ljaH3e8/3G7zDodVNJFkbxNnIRBIyt0qOnz7SBo8Bazsm
WzSKHKMTWekiJ4YkntdsWG1kHG32QUP5Tn6K6hyjbP6Z/wpDqjI5cTHSEh0i6z6D
qLIXaW+Nc4JwjSo28vSaI47yyvHPr6DIMJVZFE4/dImYKOCWRkeLdf2x16IDXvqZ
n37lrVq3GPMUq6cdOLQ9GFYFsl/54JTkA/TfE7IWNiA6jzeyy7NOetGsCK1DNRNx
r7iY7LZZht/LLrhL5+F99cy5VjC8FsciZen/VW7Ai5DpyNI2aDGAq6dDvukKf2Eq
Dtl4zx1aNebiRTbDrvRJMYxhhVF17QqZwgeZJDzm5AnzfgkGTF24hRGa1JbAouo8
PyXFp27ep+hRF+UrVSsg2yV0d+51AFWMNfmAv31JrncnIJqSRyGsboEP5FLxg0JA
58ctlUFpb2On/LJtR2d2y3aa6d6osSgjpU0AhTqIcl2uR79YepsPjrsSlsYS9r1E
N2LZbFj332eSAF0ouhaGnm7pzF8sKOQRj008eXPrnQ4ohzhrZiNyTc7Wqfe7Edzb
w3Kdo1vZRWqv7WCOt0dIbHn1Y7m76TbgYd3zjNtrnbMxtNUpWMnNJK9wm6Xx8ueV
OAG9J+UijPfptic/siyuAhIjueTckpWyVTy0jJkc74ph2AZWhCRFIOR4inTbIgzG
94ocwPEz/G+UjAj5J2ZtnXnX9nzP5cP5Uhkn7Yf1B6UwaumDnhTtpvUqnB0EAxpo
cuip9NwmCPORJJugOFF9HSf1Zy9lOZ8CpIOyLw/3rJno+sv1uTx7M3eZ9ts4FWp2
ItLJdRLhGf+jZxvP6X/JedPKGkpH7ltCYv/p8CVTqU5JUzCX0c9cJAre5apCvVXn
c8j5UmxWOCmPFLxdoYPO0Li/uquLn1WOqR07k3BTYrmfsLC5uld2b05wXl75AhXB
8nu2RL62wRq4L/c7ca7Z7hyzjRIwaf/dp4lLxeqCpF6xiavqD8psKXZVvZ2BVeI7
kgwfiC51snR9wRHTk8fTkQXzTh+B4iM73GQg0ADhCjw6hoZtDzoWDoamkEaR8iyo
UbyzDH5s4ZQ9qIqYHUfRV2Q2wML2FBpM82pYol+DGjVJgDCGQrNceHxCj+HV25KW
3ecm88FxC1QZ6A2HyW/H2nfwhN5X+C9cpA0y8PdfayNUjCIxezHi06GAsgw9+9O8
80FYvPMnSQ8Vhmmyo+36UdF2NxwquT/N9mOFfH+ISV841nqi/jrk4RonFQis0Rzs
VbpBr1S02kPOWbmu6GlhMRfUTnHD/rTH7uYJC29BV5/T0Eyb61SbdaYXWu7RZSpf
rWS2Rxi0X5YbQbdMoVsA42hIPzVo0CU3+WQ9FQct8Kyc8K05q27n/b9p11wGOtWQ
bYFCmj+PgYWmZ9hKO+X5KIsZfWxHkDL1k8u3Vz8MEGhOcb56NAYbgLqkrbMZQJrd
v2tccAQewpmqLJDL6AxspT3OXfIEK69VMODdzBN2q2bMoIjEMwKD4T11plnjGqU6
gcOh8yJBcMuIjY/nyTY7qhmtzAA0gupwmrtC+Gv11A3mgq4CmnxyYoEXgOK0L6FW
YsFOBkUVQFzYhe1z8FZhhWcjvIzXhI56cGNX/LFK2p+938VvqTJ38MTNLeXGn0mC
DJps0PAJk7t0JeNwmbm7zbe13FhgXm3c+vnS7xTAsLuN5jF+uDidf++XwCfxsG4I
oXvE1n+WvLBzcLfT6Mg+8wt2ehgCmq3d/qBL60MKny3F6V1631Lhs5rZ0kFdzS2x
PVLEn0jH1dwijwHk8lQ5hvkUigfOUqW+yvy4kAhBmAypwwuKsSXqO5nYZD2etHCO
JpPvOYv9kQMtztcI3xnXVFMCar/T6rmLGpHlCodG9UmUvuMX46/ggInfdIz/gFyJ
PDFBhalX62pK8OrO5GCx3kOjsBpLTSSeYddtBcpWi1w8EBZDnE9WOU05F79GmjkG
CcbRexU/WBJ6/MC92DKFP1ByGJWZQPTepxz9LuMaT5zVnA8DUOWL4bCIVW0RvgK3
TayoI921q9ST3u29REw55QIEw3+r4YIlYkSPHGvZMlp772fDj9pFfu6Hu/fMpcgK
R5XVzYn12UCia2vHpnneU/1PSwYPTF4RUb9r/Bz8fBhexrPhu0GbD0cL4rQS1FMj
U4FtcU+xvjNff95VvjFkbVdrN7co2se8hbS+pLnpa+ZD9shSuWvlvcdI8gqej5bO
hg3BCqNMfKXlcuGfRJdWsZopgQKfjR8O2uFnl+qF8afBb37QXzxRmN0uKfoGVpOT
+xciY0XkxwALq/o5iEuIsw4Om5VQ8LxrLj+uH8BUBxtdUKR6WvrhRpY012nxkSxV
hunQIX2WcShhoawXlvpaqOMnXEq61R/dw+s3++wuUkeM6LxRdw3wYVbpNRyDb5Qx
K3LUxYTZjxn2G4Kx7Cf6oTCG0ayxg0aZ/qTZTWMkUeZWEumczFr/RNw1wBAyyqNV
mhNfScsKrxk2nOcVJKShstNAsGhB/BVVjOqyveMxoWF4gRhdSsZS8q3/NXx2LBo3
gqYfkhxD/lQ3XyynUBEQRQQlHzO42lBhMqXCM4zULxHcMw6/QXJkzQjlP1DDe5Pz
d/5b7QmTUmUE5DuxX898XX6Jvr7mmFPXfEv5MsqHE0PM8x0dgk2mMtCTuaPEZWLW
JBFCXwN99nOBPVx/N6SS0Jd+/72HPf6b8kV1jV+wjY1xcphUtrumTJDm76gQQWXM
cr6z7TBk1xtuL30dsHVN7/ZmrJwCvAR3dErdSNHcg4QxXn7G0IE+X6VTAwnN2/b1
uPPZPrwDWCBefXnmykaVcp/AY7wKjIzNT+Py0K/bhZCc9/Lpvo/c4parDlVHKj1M
efCEumKvrJ082/zfRQuPlzuaPOFbR5DQPjFXK7gMzHBoN8bnBFD4OVbzdl7lNfCe
eUTnzHGZtQWfMX4PL9aBvnB7Lvg/asoFYH94vdteCyJpPqiIyhy27PSYKdkbzNVL
GNs5BPRKfpURoKo8uGQ68bDsh7X3XpFtlzwd+Nj+YwdgULf+hfpmtULgl+SCu2qE
XzlPCyR+a+SwcwjVs2dCtqrWbMNCPQZ21dnXTflqjV2TzQlF7bF5EfHX5UUbhoS0
ci38djDsV/eRo1w/oM/RAfVhWR13xJgPn25SUVx+bRCGQaLyY31YZrakeK+zSc1L
CiV7qOy9xpznKUQq7ZDwUtGusVAI9Weq68C7MhO71lrjzTrJmUFUFwCwdghFlirM
uhTquYtIAVDV30UtAq/kbDNfj21GTOFzpn+r6Tml3a/3YWofbgHIaBKjNelqB8CR
5i/73ZJSLg1yliftXJgjFsojMz8mzZhYu/dMLrSnmNM1bNGGD/0Ay5DIzpUzgU1K
37dPOcXCaLxzb7qB2Xylpl7y6QgzK12xjsV3o6x7KIsvALZricjCr5vxDfFKX4Z4
JEOkHvwD+8gH6qjMDqZZUABWPu68C8dd7Iw4sCcw2TPU2eC/7eAt/9JyIK7L9XyA
WLZVehMc2XlFuf1QoTHsk4ysAGp5I8+21v1d1z3+XxcZOWNVG26rB/vnV2CCmcfF
9Jqky2NVXc2J8sIF7omT0RooBtVJC30WbJFGKQh7ZV3WUhNVHwwkGVkNXCCmXgBL
HKqQL8S9xXKVRn+ywDUt47s5/7m57zgaG/Yi7xH4uwRLlAP16sYFYIJ8WUJIQlWK
k/Wd2+PQ8+BxlTWoAcY8AJNo+8u9laW61H5WHOvDVPsbbhDbdE3klCkYpmySARAZ
N/VuwoloaaqTEf8awLjq/+cC2dsgOb62snaFe+RzMACZnZAvrWQ014cynePeHC9L
meJt+Hn+VGQxdOefDzmqKu5VNGmoV6yra65VUsJvEDI5yhkv7+8pq3hXjQf30nSG
5yR1w0ZuEA45rVuKCh2gnVfSpcaA2qKWjxMvn34WE4Zf+M92QY5IIud1Lq/Zv8N1
zzz75XisSBPiHx+Ph4fziOCwDN74Z+Bt5erRPDj5d4459dudtuSEc8Z/BBUT92yK
R4pWRQaV5Ac0CwsFHnjCz/7AMABQf7L4Ck3Jmz7rNRk1UZ+og/du+l9oNEF1sSaB
T2IWSS4uAWX8/9veEUr/xltosV6lhhzBfw3Wq1zPd1XWK1tEn+sJDi9F7qTyjYE2
MmylU8JY86pc9+y6vBwLBwKQXvikYHZPA3mRlrX/V2PjRXGm8LLsnJG/A1gPVWOu
q+z3n5wyerOUHQdsUgqyuatqwe9gLR48FS2JXR4rqtRsNCVmwt5bkPU0bbaaMsrT
6UJx4dIGgr8MS29wfgNXE+Yl+zXbMCWes3kJFuo0FSTTl7gwpx7Ag5qbVo4e3du5
HK53a13Lyq7n6J0h3wNBYG6y4nD+ZPoylBBEsITvs/3jVZ3oE+4IQa8DXQGioEkI
lTbcUwl2APr24ZzXXrPDm3ZUX62kPqnTA0KP9sWprxSm8/q/foLK3Xue9bPyRWjH
c3BSufBiuPY3mlVhn0yaNgtDdwJJZCs3Mq6ZanBc8b1yRW80pVuDwE+j7GcnN4LF
OW0CyRvrXT/zOk2wkWkoU7VHrFx/ec95IgEnwXiRbheIpTtMqXAbirm6byVceoLk
5IOUScL1/0zhZMSX5a5wwUbkTDYIGppEX2aV2IMv7tViMF9qFbikeeYWLjglj0jE
6/xLjg/B9g9G2H7pAgo/xhnOWiOrrybV/7ZHPct4PsuR+esfF9R2Df+qjlH0wMAm
B9856EKAubuQYlRVOM4XlsZViR3MZ01fM/wke9HlSzWZq3akFwJJuARKuclINWEK
b3/+mR2B7W+1nIpoBBv1L1HpcSxVFuAvs11U+UhxNvZFuGvU2HW0Loj2ky2HPf5f
mgOSfYF8GugaG1yMCOeXqSpWjHnNSOEK5lSzLE8oY/QyqWFKOuamcbiOEF1uiReH
44MpaQlRCaMmhySN9glFKQ4eOocQJeMiH8f0nQjHoo3b96lALcJ1Z7062WcF9j0h
Hj/6sSt/DIb02raK3zEEhlsROgCNabLIbURWd6Z8NknRI6tzs2kwUuLUTtGekW9K
Gi8oM5fA1hdrKVPkq+57orrJnc292grnyzDjB7maFSDjBUxjTvYXBPngq8qROHVb
6A5YpzD0xE/1CQ741ZEfmJl51uT5XdfhXYqMmavBujt/gJIiOpzfPsYyuodHPhjV
PN1X6tkrqYvURxM4hKEmIsOK23V9fFyYLCj+W/KQs48ibsrvd1Xe7PYWnh7ib4yL
pf5it80GrkrxtVKnIwoDY08g9BXZPCrFITdwayewPSAZP2B89XFxxxg3GXgpTLIF
lOxakuzOqlCHAVFHWJK335Stx/HMA1/1Aethrn9eskJPpG5rG7zQKrQcCLJ+tvRK
dEALtdbOPyEm7h42HzgOPVDwNUSIiCFY0uieZHAtPqwgFHClPUW8Bb0fW5HYrtlS
VAsvHykvj10cOPesuDYgt8/2FbYsM4o3mH2vlldV0Ubn5lOGcNdfQ9f99Nel0Gcd
sxJCOmgxV9yuHbmUuQoNbGl0eKmelBFgCqPtnwpkyDe6p5GBefkQDBQk8nnKdlZf
K1pGCNdrltqX8mIyzgUc51f23velBtp/7j8ie4b+641CqLaolG9e+ETqk9wc8sY/
lZaGFawdNAGA2OEtjNa84eCHjN3zhn7CyIRfm3cWUGa3D7/afylX1HV5t0dTCYxj
cf4kzJXZaMxbKP/rEgPuBfzw04vmy1XUEzsq6UWFMnXmykR2xfbsugE9R8SAG26m
0hHI2aJDTN0CAI2Axl6PRBFujL6taNrsc5YojU/vJXsDy9iKvjTVB6IqUNSHBvXq
gPECpy2aXssSbGmqshe1IakynvTiSvhQ0Hna8KsHHulH4KY26TnV5Sl8AzvPM38p
WEXdXEiwU0l64+q0X8wl992uAHFFa+9sPZDGjtlOvR9aEEeBts4ec1O8gGzjgdVZ
xjMPbntA5a9yLcBTyuOlLu+TVllKjptP0YgH82I8uQrlhD/Kp24dS9OWcH2hcOz3
BgjzjYzmPtQkouE4w0/T9iAG16RoY+jX4GSs+yYTFxjCLW39XcKdGkV7P5aEJTqK
MkYqZ29sqt99z+lx9kcn6KKDdu0VqroL5adT4gvzaJr3i8oC+k3cenAbYVhjm0jf
+bF3nDaoNkSZgCDtLma4kyBgcp3GssEE07xII9bH6O96iJuek+j8z5yPzOUwca2z
ZfCSF4+dLfNsZgl8xK174C1VlUOO6hF5L32tzViN34Baz+fzhb5XXuaL8VNkcKnK
MBjOzH2PWWvdYHQ7X4MPCTEVTKCMVh7jELBkOiB+CjpKfztJh0mLKVyhAC+IOCDq
Ras94QVTqUddAVSHbCp/SzH9XMsZvVmaD1faEzmPWk03+ehLjSCgOsESJU5nZPbE
ZHJjyzwFSTE736Bv9Lm0An1ZGZ0dh40pUSvy2M1PoLz2PQou/RNB71z50MnViXOp
w5IrFNo1YZianHCFpgs+ffTM0z4fQjKAwO7TpfZP6LnUEnE+bD7RFiUw4TOwBM/U
WVfQOdt8zveiS+ssjls/UTc3PgjeEoGgrPOBiYOdQkcpvAKTKCkGgrehwuLFfNMu
SzW+dqbUVS4KkpNcJ0HFnCUG7vnLdNlnBSf5MT76zrWGOBFXHBgOyEAQYra/muHR
+0f/57YKUdIoo1NGdehN4bA8umXI3Y+Mdhu2+x2WFgKjWypZJJgIn2gxroTGZbkR
Nsz8XSSsgFHzmihG0Gh+tVTOnCsgusIH+sKas+4JUmxTjC6PCPhTQ5Lg6xfXrUIh
URN15l7oGP6OYX2LPyD4y4k6TNvEoLilm3kgOT++ug1IyaT2Sc9iIQt/chBTNyM5
iQ8zv74ykvsE1dhqlnarBzpbIeEiVMeg/MNDNXpA98fkN67cG9R6T5Ejhvukm1iC
F5//eEkdWXX7ORm2Zxrn4v3xXDtrx79hN0NiZnBv0py0M0Oz4zKPm+8MJBKnvZZw
k9XPVKLVd+tZ8k4Df50tvEUzc+UBM5cXreeddCFfg02fhbpyrgk5m4hV8Lp3rn/+
iockSWkNswuSGaqpz4To2oSclNmixyM8tayp8P+sMlcfnYvk9se98d+vOe415ww8
duuXYtwPRiJknTurhuLGkRjJxp+UuvXWdOJwB9HtzaANtfqRnpEf6VW2ER2gPDHm
QmeNv1EoCH2MFWShC0KG9um3diXkkkdpNd0gVXG5OAbXlyd3oghnkPrenyuheAea
Y0feEAy7DdBd/VDxYTEDgMDHGvIPzzjwk0h2eT8K+SviL0ZA9fOdE9N+kt1+4+Ky
brG2dy+jBVG7YFVcEqU5LlIGD1I4DTykjo9jBcr0FvQzYGU8ETJVZqDQAgYHc35Z
RK84K1A+0uZFWC/ycnvyAPc6GhTTAKwIvSfvmxxYhED8nZNuplz3x8Sg7Cwp7Gl8
pPiwE9eWTr/rhqdjCzvWdjycn46AzbxfmrinerIowdM9Z8JxvF4JBDdO2UpXTNo9
JNjbPTMClj6tGB3I1ctrFME820ll8f4W6uXOp8nu38tLpxfQcfkG6NwY2ZdVELTj
AK26tjDy8l4u7m69M03RBj7WX2yvCxnDKwwPfLUeqfQ5kKQp+6PogXnFjpMrFi62
vb480fy8vSPLU52CyHtVtt9aaaNtxwYHgUybkX5kxNvgKCfoLlDt44mBFSFVB74t
KlZt9wO4ShhleDciMaHarSDLmaLD+uQMbrkOUVFEXPWiZw90pYYaEClj5mZNKqNA
kQfstD5220ceQ0AJ0aDk9xU0OkSJn0MzHK39qO2Qb599kFlE3M9bCguzA6bMIhC3
IJafCa8TpZ4ZW2Ine3Qbg5MzvaTNN9U/ygyFnKu29aFSagToyc+13kOMIx5GOAto
mSBJjJerlvWotDJzAIDskFxiXmCX3/U6m9zl0hFzRs27KInfFonnB+lDO9Q0+tOb
B2h/XLQFrSTL8H8AuOV9yGLOdOFiHePyvHb2vFFAHpyEj0aYFmh6jAin/6CkD+GR
187LXk0/tTcdfyzqf4V5CZp5boq0+st/AGpsjWi+Of6cCICfGLomecjmFgUeeeGz
ir0Ipij2++cp+tOb5k3veg3p3OuGilNrFw766XRpWyjVn/AH7lEDSycOQF6NdxZo
t+y91p1p+VDSd1CkYvMyb5KungxO7j7LcMw06DfEOiKM8J53xgaHeqpU1R33uFLX
wgSaohWis4XrqS0YTLjQD/sfjOz7pSpfMVHL43vW66XBCRO315yU9Nix+dXTg4DV
FrLCrpp6Dn8NYyJdTVFaLR84ZTism6QvwAYZagDA7xhCrCS3QrYgyxq0/oW1btTg
ebp2vBeym5CWHUZeg6s6JB/RJQsKlcIdG343w9YdFzE+LHZpZl4/agEtYbq7FdQ7
MRxrIazYXXrHSh0VfkeQ+I4BK87sCaHRtHWqPOiii0VLxQoK/HaOAx1Q1dh/3+bE
LAK2RSbMHPV+83wnFoSsVj+lvnkNywc9pKqIwJMPDcG2QBkMBiYWA0KKu0+z6GLS
SAhzrKzS4B1X4eZL1VzTwvhp91cl6UZlx8pvDJA73MZSu4uuYoDWM0AgZvkNcdmh
e0N30ySggdDrvNOIuyJQdRF/Ww0PzZ0pVJg9qKi55q0JdMGPcxBBW+x58QSoh1Ul
fruOja1SJIJrf0fBnTMZDyLHxqyBy5FpZF3Hn5qsRTHaHhaWOQr0XZ7knchuOPYo
pOt6eZf4LQxUqQdrZJ1QrNPsGr+bPsXFzOhy1yQd9aT3VA5WZP4ff8krdSC5ehgx
ydBYHRBoAN/w6ctKelc5+H0QHJ8IwV/pN/XeWymz9blC/5XbHvyW9j87zrN6czi7
PfTrU5ONPgm29NmO+hP8QgzXHFcjXSUIT8dgIP4CtznW78HPe6eawee0qY7kX/hY
XsxLaxsURs7jTCNi8/XJgNBf/FTASbQU/nsV8l3ANGEM5kPtGeAhL7LsqPYpOfhY
rYAtgkjVwwMhdOIEnVl4m8IeQzQNKZFIVidP6rTzFkRHd16gdNGCCkD+Beg4tDIG
X8hLOMr+YWyWH7IUQo+q13GU4GDviFVHb32tZ3qqy1UQk8499aDikBMrwNKswJJM
XlOC+xw10P5mpKinLIi+uPUWeqPGLAubsl5OwHTdVQQpTVC+vXggEdaExTUXzScf
+xuisuJWfs+KY2Tc1Oigf+swBVDAPHM3USX4VF1b/CFd5TIKwxsFgVdmbdlKuWjI
kI1KDnxUzlfAK49cGUfXS1gRmRQgLx1RaqioivJ7NNqpv9OIG4716vRNheYhQBVD
E3VFudBrvYnAoZcYybl4up4ooipaZKt6TmMEaa7L6nNZhK6FnFTDdJTYxP0phZUd
16IY9X+XS5AhT142PF2IOebqO9ELdFuvGhdjdwiCNwrIkuulUcUCDNlNMC0h3sSs
KAleq5S1P64K3Cnc3u7b0pqbHjqr/FYwKsqtrGCon53OaCBIGvfcBxMTMRfiO8qW
oXl+Fvtv7aoKtRbfGUHGPNBgPpu3TQ1oNaVmnsRqCVahfesJDhFPEL569tF9vxfP
pIFAcfO6lpR4UBSxgcAsoEfjb84zNjhIY3X7/3tqWuMwyHhOGm1JEdApFaz7CoAL
AbrHopflP4mwLExZ6XkQhRIFLle7h72z3UeR2VRICOCVU1P+MWXYl/Ji/nV5VZNJ
cGDYiTB+RPszLBR+vH9vlcPmf57JuJeSg0F2l0uJGtG8amZWxZdOtaplceZPHhC2
UZcGkzDpiMK3QD1nfge7plOnwS5tRIUuFEMVNad0hczc4D791I8BtWV8HunoYWNK
5MOFQW2XCdZCdvBsPvWaxB1hcJK0xW2IIWKX6Whi7FNzITL+2JiifFRrhpCc+wcR
BKM0WLAfzMRfZQA/REM1cMVXWds/wy5fkSDEMA8IEfgh8Lo9KtLHRm+/1oKX76Zh
lgdaS2/eQ6YgpEKQYvXEwsPelCHUTPXWwt+BYwBSBAcE3ZWg/IxOURANKm1BfpNs
E//9NvXYg1SA1eOTITrVQrTWZmps/qAXHtKWWm/Rm9a0QwZBpSx4ExY2ZRb92VfW
TyhmZ9YpTbDBWz3DBqEbWh1DEETbZIHzhIMR8PPloiHq/LZQ+fCm9gvv25w3FwIl
w+CdQQzrDvBB8sYp2Ct6Q58Bh7PmJ9arb7qgutgFilJ1KLhodTacwPhF2ESxA4ZK
fZpJzOPlWN5xzbvWyBZseuk7VFCmZ4BvPr6kS4i3mnvMZf/zBIkXVYQpdzmPR08x
vUoLhk7zUFDU5/5PLUva+HRCSNANwDHsKn/4en1TtAoGOBBw3SU9eCkUNpV1oJqJ
FFhoUgFEe9dRk+gEMEIDwOF0/+8ndc0tTKgAlx+KAojUWJZMKXAOiTc6/QbAIXQ0
Nsl4p1qyyCg9Dj4vSyVAjDzoMQhfg9cp0Rqj2DDzCQDpiEKY8NmWVuX4s9F+2LKe
1iDjLhl3gc8WkkNbCsunKeHoyRjtLaJoI3O97EX+fwa5uhB1STF7ZfpbjciAA1zO
doH63FvbPOiSg2+VaprQF3H6XxtYic0RfP72/8MbHSZ4i8VDbkOabhxGwytzjEei
BmQ6XyGDw3otMrmhufU9zUmz3BEVRXQc+mjEyyU1o2mrQZp9zRRuKIcAJPVHS3dY
2gseaeeeHxuZQpIATvCjLN9HLiCRHgj1U3tD0qrEfzNKGkIVmhuGATIF2kpv4kvD
eoeKbeH6l3GdOGIngA8ZJ5Co0EOz+aNtvHNJr1BNIvp3gXdtZ74G7ZwH2N9gfYXY
eb7VmZ5ujyCgXzlewCx90/tMfRLEFqTssJ6cPctIZ/Fux5jmM0chLk6+8ROyUXBB
PgXzc/aQcAufgi31cZnbdpzCUdJ9DvLAIzjtSVv1EWqkepqXu1nzrfPJ1mJTLvE8
9BZMNRJ0iCQN7W2X+GFU1oR5f4nvz2NnSOz8e0e7nHiyVgyBNHD9fvx/kUwAHrJE
AEYOoMAYxzO7KWibZ62zywRacFkV4Qba0B4HwrfNdW1sZO4hMM5z1EMatTk2QpsD
Fvp5M2dJk5fm9ao6F0PWLFilk5R6nLZENynzZebVxUyO4pKjTX9oZaGOImf2zH60
FCjS30L9q3NDgD4lgaP635gJSpId5z5/2FTgZDEO77u2KBoX9Qk7Rdkuy2A50y+w
wynl+1Lar/GtDbxyLUWN2x9m8+woxbgN1Lyu0Ycza+McIznj56WxI/WwECI8Qmk4
azM/W3Ab80Jng4H2FJ4FAFMswrzV55XHW8/t2dEQbPLnUNPX6q6JF1iXiXFgzeTQ
Kp8Up13UwMZgB9ww7Lv70sTQRgEEAQ3/KBTU3skTBClyZre2PihFhZt2vDlrzU7b
d5Gqo6mF0GiVC8EG3Z4waKElW457U4Oiug0qdFNsXx7tIEwKOA7k7aWF4w03yCc4
TbwSziCRwsK6h9a42uZSEx7y9wq6IwKgrn4MDB/9l0k6H9glnCNv8EZo9mbKbJly
qpfvJNSzzn0+HexZXnzc+NdVBpF940fH0UVNS+/Hzr0WxQE1CUlWWY2fUD82JPYB
oI9pMY8WWbn15pmz84lDXCZQ7LeTdpSCQYRQJsxSfEaITZ7kXYKcvEhJVGdcK0VJ
Om+4mnSB7aCOMhGYFyDugprzz9mXsFosj01SeG8v0DqvJotGdtTwdAeLHhXJRWfW
M3d6AnQGXqcpc6gXip2wJ11BbpkYyf8cSqJ9gu1xuNLqvA0MzQtE8QKaGDj0tqMV
tRLYYZ47FpJV9iM9bskNiQkXprS/B6VMn/wtcCmNrz4HvDREeCNh9pQAG6Hne2lV
nP91fHZpG4gGMVOfzBNerDDeBB83h9ssv5/Z+3embCW7WUMGgOMWxQNhq6LcpPui
QynMvO9NZHnM+v1Q4xo6edHQOnEfMJ1jjOe3bOX064hVDq2Gnxsegvdbb4nA6oX+
62wzVtTn/MXfqSBnijWwlaNd7juaWIgt1fbd+NUYS/EWeX8AUpxZRveSb+pMhzbj
DCb1b5p/WOe9F7DCEKCk1ilofFnveDDjor7u2kp5vcRW8cHwEI52PAPfQJb17cuU
iU3axA9x5EQhmzrRIPX9i8AX7owCXaE9O/4O6Gq/AgUMbqX+wc1lhjxD16LL3e/U
+VYSenK9zavKKtWO+fl3Lv3UbNZ+0lwXwYTfB9Yunh/XSjzt+Bb976DQlYJW7oU2
o/KbGRoHsdR1lXqaCAMO3AMRmHwst7j4/uygctimR5KF9am85dEjfmPEGZ771Xen
SVd2zdl2OjP5iHiJLkIPHI46KnmgytfKdBp2NVZKbXBUlgQYpEbKyBYIFK2vAKpI
Rzo6u3eQ/8VC9d6tB8GdGed9EKNXFw2zarhGGXTq2TKQgiClXmQ9q+E43QtsO3S5
+w/xUWxvoq3ETHhCBVJrhlDduaLuefnC5NjGIJCOD1afdcHSsb8YaWDweIKV4Vmd
CBzSeJbfk09rP5i83azQ5j3yGtyxs4mDVGJvZdQHDVOCwafRsBS3fLOu+Ay2h7J2
YJN/DtKRZaWph5GAbu4LlzQFGPS/kyX5fEN61i5zrFj+YRm4o04VYI9pDvTCK/ej
aBs+pcExDzDO1QXnjOITMcNqGVN8kiLI6dPLKQxTrUGhrdh8vhFzzR0rhIwjF8KZ
Dp6X+EpXeMLo6P36KFyr6LoiTZuKLfI2JInDihHXij2fR1oW4b/mjuR6n9XVqkV3
ZGuxNWHyhAPvl4l68cCPjw2n10ohoJCma4se1IKsLzZVUmqRYTWeOreep/ug9z9X
UAShbn8QuWG+nducLWhT8CZ8eYYPznRXRMrivsju40GDtfi6NFa8C/xuXp8Tdth8
cmJ2tccnVrLgxqeU2A0xuRSPP0lFC5jLASto28dXg765MDmAQ5e9oqcEgHZ79VKs
OdzGE6b4tfFmfhg6mshlKs+6GfeJBMSHWsSdunfz003gF7aT9rYauK7cqQkzYzIQ
7ymMjtkqN9XT6ewcP1mM6KM05rUyF3Hq+CAZ+6iF51vGxMMQBxRuqemL7BtA7uGb
TVJawtAMJucztzJNrk0j6rWEekJjpgSys4nch4S2fe5R+rSaQogmQURuFZOY3noJ
qCYCa547oKFeIdScSR/RAPuOvxYK9Q1QpWKkVsLEAsELTzQnZCYmtPkt2FoCbw8N
AO8u10x/nKXljmPWjORkmPPJF49APFpwA0+F1YDJcdCNutUuCGowLMbHPuMQ+XiH
i0FNKdW3/Gv1vrXJBU+5TFaWaV/5WNKUJdecP1U1IIT7XpsM0PNYsJe+cpnEArxw
SoOjMUeOBlkmh7vRD22NrDxwUKAcMOZNCCcyv5KXh9lBi4oMNxafuo8TpGq1gJte
n8JYPgq9hB/RSc6UXRQCCLSsSQboyP+OIS9I/zjap/pyV7OZNnFv3qLGhDTxCpvZ
0k9VVG38Ri7or5IJpeLWicXY1+3xAvTEW0torLiqYj0pMO41QPiMR2CYH9/rNaNG
Fwh89u9J1E01g5csVgK6M+wnrwdqfWhSyvLPNaghSGqxBPnKzIzKJkGOsG/Ktj49
x/lqiXEyyHZFEpC4CKrA1LcBNqskccQdzH+EmUgygnXudmPI0jkmDa/Z0bbuNgRZ
Q0mh3LAkNR0qwGar6bVnAYCQPFCNvIVCDWZgQs1+dRsEIelui9VpTE+1+Gq+TvWF
S5gJWt7t2b83O3lcrm+lh+AzquNPz6RpBNX3mXi2hHSz9TsLqMDpfwA1hlgb+Q/V
djWhZzDz4Lkd2AJE/wY+L9q34VEAAYTIr9CRaK+YdmDEdfU+dvmYUjYwcxnh/rOY
Qm/qRsBXS7Fykk38O30SvLqjxHOFRUsaaEN8Mp4cn5S8lAOvFTUkFKipmx0oxL9O
9+rDReUN7XeW9LRc4t8LzqpoDy1p/bfXLhIY8wBk+0V2Akxk/Tg1HoQwgdw9Ozpa
EU+PaHFI5IoWa5m4YYft/GAmviHmg1Pe+UMM8hw2U/jnkzn5SfQpFvG4zsQE0rSF
68o5pYWU0awiQ1F1mohqi0l38ND7pH+cNetiS4kwmMo/5Hi5daesUhe851M1z6Vr
4T1rFOHlDLU7a2tzjAYq6iHpNplWnY8WYmH/dEnE0chis5jx4ymO+g0KL6/i53QV
cF16dyd8ybKWOu2BUJdO5n5x3CLO6ZpkKvxKX5ve8pVB9ob5NcJDpqMlaKLMaswv
FXDe3EGarbqaQkedQsAaG8ou/rT2fuyzNuGg6eFLS6wZCjnpxrfDBM8a97YacjcX
tgR2QKjL+RPo2fIeQxO+xlwA2r7AMD9oGRsrqkklKMUPXpKzr8vSynjaogxvgU6l
I5nGwQ/1wvuRqF26IQ8DDgINY+d/h/14jH7MhlrScQKc9ptnehwf/2OOBnCmlA1+
V+DUpK4nDprMonvjbuTPLkuVeDFqgrPGghAXVXf2jSTPjII4UBDCIPpL8IfJB3uI
9y1un7oZkO3VAUUD/ZMWZmKqC0vgLLfEh24XKkoL1dYZTJs/qML6eL9INv5ZI0JD
+WF/VrIzwzw/frn8+Xj/TnT3MQbYugMT040H039iTZ43IoC4A0YiqRntjd7ATUvf
a9gJVY4AwHEqEO19osrAZE+La5y/euB2/7heUJKUbVH54ElhJ/QypLa6dEGgIb1v
7EE41P309czAOiS+XW/biY0Xh7DLwEyy9/YDjejLziXXuTUPKf1mJp8xGMy3+9K4
B0U5Xg6n+1ad7S5dc/sWq9kZ1gc+vqmPP4B2E+xV6Q4Qhe+XPDoSm1JP2Ymvf0d2
79nmPuG/c0DApMYbHjQiUYKuSs45ji2qdtbCoGqvSlkm6hG3N66nmzjvVRCvJ6dr
ZAcHjZnEDyuFiRhQaAPZI6CTdixHzS74+xOfwKzNZHEETl7ZeBQfudvY7EsooQ5M
i9LiN3rGpSgbvStFmPBuVFqYtMYj6kwE3ql9aO0YwBAsL4OnWMr2EI77b7V/qycA
zQnu5Heu88r2ByHSK7qfGMo7BlynHCJrs7jzr7o8JZ52Ybh3NipYmGaKdVDTbERQ
AqlzDl88t0qrvZoPQcv2dXRqcYb0GWaqoOK7eI2F+U4XTWjBku9p8cM8kirrCV4n
F5gouRXCtxZFuIAf0G1GdeBSjrIDrUauuZ/gzibwlezSMnGaFp7qKLC4QMiMfusA
wADcXZ18lN2TJgUobPGubE76AjjqRQh+C1zou+w2hvq6YMNAgBOGrZeYA7G8bnOw
M8RU5tCft0b9SBUusJ3AxOleh3YLw9xY9/WVI+clO9VvDZNFbPsxjzr5KscFzoav
lZEUMdkXdsaYmXFgoiOME6/xQFvkJQGYCzrfj4jH+1yb9DBfpWYLFieJQHjhvUNY
zkV7vAAGZu+LiZj8n6YZEZY2Z3fAYMsH2xqE1RY6GQjR/1UIlvJCDzpdBgcMfkBY
gu2Dyo5rV5QhoT02cd9GVpISTPdNH6KxAb+Ukdm7rChOY+c0Y1II1001+YnmIU1M
Y1agn1mbw6Bbariwlf9bUBbA/dlxGlwVajRidiB0DtlZHDfK/JZkvXidYGJ3KPrF
Zhsr8r62uAQr1CyBxGnO+ZnbMIJ/Uxt8Qcck54eLcJC73/300RCsopRh4iPPor/H
80dC8eEJDjlu/9VpikdMH8V2dbGWhEc9Q4fn21/PbKzaScTldV5OYTPg2WUxvYwr
x50JfAOUlDh4BKtrkQ3hD+eZMo4n+Xc2eSIW9lYGIQG9qLAsE4q4CfYvKQQ5r7G6
5Yq6WmT55LjsTRY+HcyFPg==
`pragma protect end_protected
