// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:38 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
psYz0ZlGv0mvmHaTAdRy1R4CdMTLZR3nB8qBzoDTYB2R2xBsurUxfqcVfDWmQ68+
XA8BXbv2Stfwdcz7pWAHZp1dnpnFjC/THmBZhI36TjlsJeTJiN0ZTnh/qWOXzLAe
RF0z48xhko6JKzZcSwKzLoTh45nWZe7UWizFpw0MD4E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19952)
rjBuJYhHimDTGCExvlPPx4kxSHtiaUIGzYcycQW/yc8XygeBdODZKMu0YcUxCItq
ijRJdULjw6xjwv8pvnUymUm5tx9r3Aptb2vssLjid1pC0V/I3hfLwLuL9KctJDK9
tHuUkvY5KhH8xHHd+5sY2WHEFKvWUjxpOemL/9z1/pfo8KsRr+s15CuiOjv27dCf
35z5mxxHaKyPSLpy/ctO0WBTsp9iAx92ZzR+UzFkLLlGGIXy6cqY3duQWqiSLMuL
HY1Lwd+ncYW8MMSBWmIYBs36ix/vGwwMX5kKsonNRLtEaP5fdFk8ka51qwEHBbiv
fC7FJswvx0GzhnIL79kffTJ7bY4jTMKPSbFB2YINJVsdOZswgp3eKdXgYxFrA4kf
VExSLuQfBbY9UBgC6IdiSoWK5J4qR0bXvD53rcKcLC65cszhYBiFN4OGsN7jx1j2
gpfYt5VtBu1XKnEZM1T+Dn8G9d512hPIcgfnX66wAGTXJ/f4584RgHgq93mZw8fx
uYVSte5w5MWPzrGKJkdIMVKSjues9P35FwTPHt7qtXkMETgD30yaDwCHiEn9sh3R
R+wVe1p3S00gF46/F1l8STTRCBJhXOzBb7L+9LqI73JtNM0KAR5kqroPNdKvC6K7
sbVhnYbt1mJToNfqJ8/5/0eH23NDxaj3qiRtnDbZCM9Usik08glcCHbHRBQ3tu4N
Mkgj6uzTfEySNP8kI5fYNABjdHmZvKm7Bq6LX5GZLRLMWlJu6Fpdi9OzsmUKkPJ+
e+/8r3giMDqw8NQyi+Xko61eQfuQflI6CEsj432hD7miNeXm9VGBfrlx9RdviO3I
PCXbHk1dhQLu5MjAM71GfvGdWPb6b5J34NLpGPDFkgrKdQfB/Oc1BKMwnZcxvViw
CIDhaLpx6FZhLXnZrO37qmoMryKJjNdD+0Kpe24KqJZF0ZSlmpcqoxUIJ73RNc3M
dolSr+mAtXNDRVmgZ3WwyfIEcuf6aQ2uDTwgeeMsYrfQbWLG3PxMLBr48cwuqCtc
Q2b5cRdIxTAd1dq+BpFqEgCWJjc8UsZdO+gxISAWI4U0C4r1lNq/rA0P01/ueuXv
LiIoaBCRxCZ6VdcZd4mPdjQ319w+O81hNkhmcbeDO8nJ2rs19wtYMTf4UxwZ3aKO
ceR1dhZlPtGtFcn1vVANrtE3LsJU/vuYPUBPK92PdFnFwcNOE1544VXkzbP6M/u1
9heoN75ipF8tzGHmS3EBosQTRcA6FWT3mt8HWoeGXZiUcuLFYjS6i+pgxAWF321Z
bzN8aD4YWy5tgDd8vphfTbrdfrHqA11+g7UO2xEFTwLmf4W/mNKF3MB7CSnTV0cL
yzws1sD+VwUQyt+UVVx/gDpn4qruEGduCQi5My8hG678GN+Vc1NLRGVqHuSrAm3i
AVzmj05dSldXVhUyRIhCRu2ZhL77blP8NT9fNNIKKeB1xr7MS5pC2BDtgnSj2A3j
UBIAPQAuXycQcmOsh6QiZHvgfA9JiMpqoexZ75w0zaRz/NQFfH9WWxGQLX5YvpdL
jywuU4mmFKwY7unbZyS9W+VoSv3LQI56RHH+wlqXZGSx+UgoFRbfaRlYL2gub03S
M0IUidC1BADdksk67hu2gEd9k2JPU5G2UjKONbf6gj7h07Dt8ruDk7HVRHBbjcq3
AJibjYUsU+dk2ptuRWrPhJ7cRXG2XOh1hYsVlmfE6FEDAEkQfzu6wBN/1jIgD/m5
DRHhM9Qng8o9xqTHX9cwzPOo4rSJWJszh9K570xquU2mjy0NLA9HkA0ZhLGjYeuX
Ex1Zzc+5pOfkW6HJsvwxG3XIe+gPJkjJt01SMBiTP4/jKudwUyZSV0gcOni8JYED
07fWOjvCxTU87IFfyKggUFpS/ltVgt2KtMumT9Yt92+J+VMP2nxtyrUfaia+l46K
drLb6v1U3YhbdIthBIXFgBq2k/oCynay85d+PXpdGAZHzE/J5uVAC3zh52/vjsoI
itPQnyXXyPWqnA1+RyeobGd5dEwSWj0c4HV8Hi+sFfdnUGAWwEu25oqtZVoJ+uk2
1y0XMk302pRCTeJ2ZPHf4MHNKr7C7TAC1u9MK5U8uHpwrZGkupsmIXUTj3Gulg02
e5Mtti/LW7vFOOmvGJ06Jn9aDiftp2XTdV55ldKtsE1zKvcWFwiXIelIIHY3ON4+
1Tz85mLTd139Qp6JG56HJzH03ruU6dNl02GDUZAWnefqmuJcpGS1XPI11UQO8Jzf
BadLWDAD4wRMV3/vWw0rsS0bpQrYu99D85bGpL4fqudJ1exJxSyoMQQZHktiDNMQ
gH9DjE2ZWFEKqyLM2+fyjgYY3X5SltuYcQCB0txAnKX0BQtfiaXVi6usTveAlTYc
UXIgvd2qeZoSaePB5BgVFMEHixuqIJFFnlJdCwPiYSZ1v7/6GIa9gPCvrkRUlRcF
TbBaNOS/pxxfchBjSDrtjI3K7bxOan868ao4alfS++5SJQ2l0+3FoQ9W0OXkbNXV
uqciHguWuzUIqsyFym60Wc/F/3KuF4ZWWnDp/eu+eFf/EA5vDKJvr3x1x5jeU09t
ZgcSe/2id9LUMQMCqFkCwoy0/HFQeknPkUd5qzQ9wx0DSLvhStENfk/YLRJKPA2f
5KiCq71OTg9aMYutzu+Nwb1hjaGNBf38I930GqsW+nKbikW7TpP20fyRjJYWBCM5
ZJTGXdcl08Ipt6lRUhhCuU3/RmvZ+3jHRyh46LESrzxiLfeED8jWFwm2XjI8V//9
MsbQIcIY0bHFxSauh+9jNr9hBzG3x9qRRA1XViKw3W2i78PVfTVC1AgUGz/S0tBR
KjeC2t/DOZ0RUtWMEu3zkeADMNEwxS4nCku4fPPbwnF5jfCrGDb4rMNGhKGXkmXZ
gmZphLJge3iICyIf/YmVWmMe1DK+55gAH2uRKUkCATvv75it7lQ5nQGfmWVqTmtf
cCwli+JLbXBKL/vcyz8J6YEMNQRwlQI0DagZDvKeIj6OpqXamc3hwhmjIRG39BRv
OoSORYoIsI9gCynCYgJtRK0lJe1PdSoIjWGm5jkm3AtUWiQnYbkrg8fDx92vWMCz
Fp63lkDey3CK4F4jR48fqwGToseLKXmAlJ4SLUiKDAlVtgkVNc+hZnaJoUCd6eHo
YkZaMxsfqq68CYmnhvOq1FxU5Xn6J2Yrf9KuSWxJ7H80nYeyn3ZHjfi/KvPNmswq
sg/mH8ZGyJdc7fz+FUDBcybbTwC7S0HK+mTWxz3bmrOij4jDoGO52rkCFqzxuYyj
+8ejFYV2HyX+7ZE6viIdmFVS+NiD/LfP1ahG4CEvnvLg/cALey9uec+UH76p+MM8
P+N4lJC2dXLDfeiw9T04c0B+QoM5vus/TdbxMaCgc3oHpw7FIXtWUSRJsAqHXoWw
Q/pYA9bTgJBeOW26ThcTvN0nqyeE0yWxCxx+QvwFZ1Hf4BWWSM7Pbv4kuxL+Fivo
m2zbWVTj6DtcF8W+FwqvcZJVsVkTygR5ifBTBZdtlTikzV3J+Col6tnwgLXa0zgG
Jj5eY+GrVDUria64WfGxGQu9bVkmGlTdgyTc91TgqKKx6+MCUDlOnbXONee0V3t+
vWylfElZZgzfQnauM/khHxwB+uJWm7K+V9xusqzT7Hk3+j6RKeJnbrShy7qHzKtA
U/FoBiUOlWCdKUg9dyJvHPwlbOUzMTvrna7yBQWY1qWTPA7zu8r2RlbffK5LAeVF
RqqIcoGRJmbAaP2Nr1Vx0AX8SHjXnGfrJxI7ggp5ALpuFdTbUsl8M+37/CJMEqXp
fGovqqEyteIUmeJ/oIeJguawZaE932y+4kBlMQRF5OmcwBXAaLvMwKhQBqaKiLeQ
87Ch0eHfCUfzFrNiBLUiY1hCY7IQ0ZCQvun8pZV1uYr06xBSVALkpy0/4c6PKqcQ
4sx0Z7zGlikZldcJ7uGfFr/4IHqoSr/B4GMU43MVoRuSO7Nip08AbvohxrslzpQV
X1y4OCVNq3p9QA4PoNQilgrUEuSGvjkTidy2fWFnvhH4ALmFlRF2bgtxjE7YfndQ
DNcRmp61wZGb9thtrz9d5mJ/r3hLVMJJEXfaGjUL/6NO6qyvtH4PZzOmAk0Bcgd1
zvvRhJUmAlShXmbEKdEmNRTUZuBcA9L8bjl5ASmWVlWX2PT0iUbkOGMTtqXgJ+sj
n1bhRkQQLVSncRnbSAEuIiehtw5OVuNuclXnFju/6Vbag7IhW6gpaf3wPKa9alqg
DcJhjYpT28o0BHlaTlk+8ODH6aa7ha2qSQxoypcfgtqicJc3RkegUZ2rz13boXlW
N+aptJjuwHGX1s8JNaFk5MxxN3o/DrGUvhvm8HPPmhogv0emVwzFMVmDMgsx3UY3
bKargMPj+T+wlzML/Q1jgZV77nnwKOJTM/KsTHg+J9JrsAXeMwBIfaosYAsH5+Oj
CNAWd4b34HSx1Jq/tH8d/KZ+MY4NXiTbpCT5KwnVKeBUUAZlYfQ94Y3gpPYIcWyj
K6WzutlN9pDH9g6haY7ha+UK9DOZ8C7CgtNkS7H2Xro/K/TPdBKXCg8Ex4rc+XRS
rCaN+ryN/T67SpldE4j5NpBZltF34sSFwbKiOaRqy/EugFf97utRZ/8eRO8ifqtj
CC3sebNrdJS8pBKpaKT21qMuMEoilLDRcC2Bct17MJyJZFmwpD6ron9XzYVMANal
3aUvVOPJYnHv/cutJRWhD5Vwkko5PoBLUmsvpOhDirxrOX2xD4RGa99fBWH5eqxB
2W1k8no5of+Wqgeqd752ejSM0+XC7ietbfa+r3vQlZP6ttbB6nWrsoCFV0SOVws4
P72Kkg1D2by7NkK/rQAPuklENM+AJNKz1u8OVqvD1LNoID1z7FpVXlzwDoKDnuoA
D2eGp8nub4wFh7/wq6oiLKBsVYodpJtt3yUfNuvLsmyo/Cz8Hw39YRh5crBIa5qE
z+mHhUpodxiLlqsL95bB/9+izKUukTb5esNj/7JJ0AGe0P6jVBfnOD+k8N+VV69g
YyD+2sbWDnYjsG5qFfoSbMJp1o2OnegO6xvBbaK0qPAyqnA/fQud0MyqaSILpAHN
m3hq8FDU1AjIwXA6VjQ5Nv4u9ZqAO7nbbU9Fz9FA52uZ3WMqYjJgEhs7wgZH7qCe
sSuvEpl9T2obIRc4WfMKuuZ6ax3aj5etjT2apa32/jdWhnJnE5vb9gM87M5CfDCb
VttFfWV82ylLzEK2cyBLF8rVzRYO+f+1hzwQuxbtLSNWcWzznEZ4e0mgfY0loUGZ
NctFfIyjPe3tfbBh+N5CLAzSkPSdIcz+tbTQkPUk7SLdLM+AqqvohL27e+YXSeoF
FkCGzx5G2lMjpfR4ZYaxymRGkKX7Sbfyvb51WUmksC+dK7lTW/i+wDktdjiMNiB0
nP7Axh3TBiPIW8pLsREG1RjrkwVwb+++9oskV/svMFCKBbphisS1cQ/kWPsietPh
q5XCD7v7owVENyPFNAt17Lb2j6JCrknnH2Y9if53eKP3ylpmHcGzLMo69q6FaVMl
JpueUAr3cNiZZjzPSX0/KWPyyzq49g8JcZ0v0LEjo9IdY7swYyiSQQUnpfaBvvU0
40jNYuMM7k4RVOVoIyjadrPiznM9qhsirqON52sE4B4jtgnWLmXpTDvyFbPIIpxj
EteZT34mCunbIGXXFN0jnTSfZs1+zcS13fenf9aqV0huEAFljFmbp+jFZicmsYdI
dWvz8vtudwSXAPCxiDoAGG5039McWo4gLxWuugx/f9Me5bwaRBmhkiT7wpOd2GYt
DJnInVZ21on5gXzfLhrNJBxxGfKjtrfWEhjoiP7JUeDPhKMM4XyxsuKECP/Wj/yb
MX+mpbVjgxuqJuUTxQHWE6Uxts8F63Jo76Ofdgzh/dNNUjBuDCZN9oUY9yMNy3cy
8TP9rVZ2wUHKiZCst20LwRUHKZ8X6eI23XfVCkZIzF1cA6Bh7EZ3feCcwVKpv7Tn
G02z0X0svTILSISTgEy3PQj0fuAvUNZrEysUKRPk6HqRK1Zp9AG3hlaYuwx78spT
K7STR7COAPZeQHXye8b25zl4rcDO02hAT27Jrfwgx1puz7k8l0LfmOQp0uXd6R63
Pszp5I2mB+Lx8tUJbgbZThyOpCIj6ahU44/aqcBEz9hZeIy5GYjtClQaJUNCCwjD
iUZi1x89708ETLGlUbZjNJPy6guwbKzYYdgTKosMZAn5qbmt+K1/tzdvlvT2SDpu
I1YWE516vS5lPZlwuCUmZSgOLojyZa1NAiFwjO5DQA5SGrGQjwZHRJwoXgTxqm3h
aA9kHhiqld89nrxM4pb2RoLTenV44XZMlz/p8vWmXYs1N5sELAhvTPE2khwuLIWs
Pw/zt3eizo0KuK0ADDtLFBI2+8gbaU5jyL0x6d7P4zU/qZmZRQsk5iipJHk3s5hi
W8yuvAaYLO47WXOZTydYeuZX8Jraiw8MQEaZtY/M2tFUgiLPNVKLgSjtyWZA1Bdy
T6+BPxegyDEFcjEf0hQWQcqholwsJGEgyUfH/vY+eGZaLX5SG2mkas5tATYMCnGD
eTgEjkb3Z9oye6ARpyqBM+GstMc/jYCyVOr255kdJP311eHKRH88QMFf+2TyUAkG
Q71Au7g5Kyxco9Lk6H+1avCzgX+SxZtuTMbRiZ/FFtQxV5tslpEcFoJpvg/a260D
7DU3zPc82jeZ6mVbm53L+iON8jZcyB9oD4VrzS9bmUPputCP0mdu7FuP9PqKzW6O
m/7OtDa3aPPqipeNNUdUOPsyBCGGkBPW1OcOLZM5Ao8ILFQ2So9tQGzSooyRknhW
L/GswblKN3pkgiDNKLrCRDefVinQRxUUD53pKrlvFPJSAirofbHj36KQfqG623a4
l3+wvskZjb+o9egkuBZeEXd4jFL845r7dLdU7ktKUhX8xUdrlBll9sNI3T5MKjWS
L3cLoTXifTmLQlep31HyOJbzPnc1pAru+dBDkh0Uuv4S/HQmSGkOUxPPpCkvj9LK
b9ZFOobl+4RMB3EnotVBJ6+9H8PHCOVVXIdOQO1EX37ZctgmMnL7fPvBk5oSFrqo
43EiPWstxVYSvWsyWUkxJaHS+D8YtFDiltdCL2corvx21DHiFvD2+bQOcssxIq4j
yCvvki00jPtbxAgWHn+qa/Otf+f5MNO35rnqpFxtv9ItuH2J0OeBul2XQGg5j1Ff
Rb5xjeRdyhGTd8MZARJYHzH24+VIADj688MKnDG6iPDM1nVkTcsPxC8i3zo1fRuQ
scYToLmkyxJFjziREEcSKeYmNdoDlmlOB/Y7X4vmFh0FAujqoNEth9eNywWX80gT
7zOxoaIbdpt1Wn+/H7WWr5rrPKs+vFxCbfXGwz+oLszQIrhxntRkU1FnDiFX7b0j
AJeyN9kqvQ6In1+97DQI+47n7yAgYLvHQs0lPByBQNq9BVCAmSo65bIm8+Zy+ZF+
OBoSceVeD+vgZxVTRSiaGVQjTVORgMFGaZmBplru84+vPcbkmwizlKgeG/nBZKbX
6+lJL+PAyYN6D9HTB5E+MXet3vR6Np10M4YKzivvz/nPLsOtzfKdz5BqyyCYUy91
jGT2zq6H75fZIFLfyDFBHV1/9DSObAHSLomeczXFyoNbuWLR28STGxgFzveoyk4F
c38meH0T3BRcI5RL7Z1dQfco78ymuo2L/s6HfWL8KaMFzu/nKLWsh2+Nbny1WXmY
qBgruyebL2hB8JDCJZqxMip+KOdPusCt8y9t6MDJtPYZB080SENdbP81G2aK4RVt
tG7lzbTel5+jS9eQBMbwCisdctdZL8Isr3P7l1VcSF2eTRIIZJANZfOAp0Io4StH
GUwlgRZjneURNuvYMLQpTb/xTBrwCYJZ/rSe9TXRbGBETKbNyCEOM07BK7IYPCTx
HTFeDggEpHZYewp7U7iLhr1U1ZLESvfNh6xzDh8Xd7eDd8EMCNMb14D137C+WUL6
hC7y39sfARqGRI0+M6vd6DcUcYIdppKkMZWriImoomsyYYuoSnEJQC1btya6mUAv
maelvXEqI58Xd50TW/f5WjqR8niLekucofcVHmLJ+0j3lcNCP71RKnXj7Q/nDZxQ
Y81jVUksh4bgyMUzyQr9ebjxQ+Kf37SJSjyiOaYZIM0jgFBnK+smr9P1YGBuhwt2
VhVMT3QZpSux04x8HepflXPUKRiIFYDHNhYkP1BMgrCoivLUWh8YNhATGMxdm+iI
20W5WFa8ElUaw7VXsHN7zbSiIvB9U18csGN6+ZKfGQrNNfvb0vrsrP3zKlUIsW9T
FDRzdBwtUPP37TtRqIc1qhLvgwSlILTb5o0/n5YY4ufe1FcyigUs/Z3y4BT+zolw
lbMF7Nbikb9IWcAoWxLCJNDD3gpYVZs0mpt3Bc7/QNwLSXj4+wxsYWz0hzTP/qO7
LA2I8O5YHDpbiy1jlpDwwaGVGm8oGJF5QRxC6OQCdyiTCLHUj/O7i4fzdsGEmYd3
8fGEoY1J4L6vgWjeW+wCxduqLlkAoVjtY2eWbx/aPdAqwi+0S8F3OYcvqcteBjN7
7ZkgkPPkXJoEINsi5tN/gaX/AqAeShhF4wRHoc4utJ1FuwvZTD9BkLI21YGnMisb
NXG6oPIvNNwiycyw0Odkv+MQmO8+UZfOyez/b9FO2w54HBTvf8br0ujX20wum7BI
0fwOw5/vMXjeK1w6nb7AxTLmtrQr5vFCCjz90K8/Zygb7cpB4Y+S8gtwn7QIyq19
6A2fiej0+wOYhzK4aVoSGQzCIwV+bIm6q/B9aUvtwggJggM+RG5qVqE0D23WNGDI
ya8vI2cVUa+AZON6NAJDNzWGLo116jokrynw/XEjANkFTpoi2NXzb4+eo5I2qzza
+CBTDHNuuCSjdueLk4p2qgIdfax9uURYRooPhcnViYZuKN7ej0h2p5uKmZEhSndf
qR4ibqhKVMcqGB8XAs8m4Rh7qiCDF6lHMNHt2DJ/3vYLN5BIUkGRlxZ0zfcOa5Bp
5CT7tJSeFXeu1W7aFRaSpYGwnZRTDKNBIZgJtfKg6KzRwaSwDh85QnuSsLyxG8i/
/wN1gKfdRbbUa7Ly1T0cnkq+0ikVy6CrdTyxCjPe5N3ylYnmfAOwi1raHFHathGL
wNmupT+F/eZu3PtDjAwxoYUQdYFoWXDeq+gLijWTKj7aSvfPUQ5J24Em27S8OAbO
3KBa5/xi7G0Md4ODMe9EVH7H6l9TjJskFs8R9KzNQsiy0tO8h7WlXKIG+O0aZJaO
uBJSQac4V8JkeEms+414hQQxRgyAuh9d3CAuniO2t4U9bsUx+oAEbPOQIkIS8B1n
FPrbU9LO1mwUuBIEj6Jz67J43t3LsMbZpqYDY1qaDCWtcewpuvl3fJrwoIL7TXi0
we6QG4KZTYGUvKQVKez3fACT7t+heAWWMLAGlGYYdJ0Paur6+omYwqx/ER9WIEaz
etW1Jy4lG5HuiXtsYSxdKPJEcsn6FuBCDR7yux46QXnyqYucjgYrjh2kVbC6Yluc
6SlOxwXPV04tiYJzlnDu2av/8FU9KVXa/h6LlkUdkykKKgu7uRWJgtxLrx9WOJgk
/TBUfF5EMEF+nGXcQ3Uf8Bw5aMTamvDvHvRlIciI2kqLcRh3vf9jmPtYHPGgPfPC
0es6ZwdzXbFsIom+H/apGQ0G7QVrKl8zRwgpFnmmy0lc3EJaOQXlZjJqTumWC0PF
x78xjZ0Y7X2uemUupDTL5gHBBKoEZUOUCt537PZy9GkHqdVQT4SiKBzdrllNyFwv
nH6oE62gCvWdXJl8rIxUrpawCgLiWH35VjLH9OxDJ9/yrt1DeWenCel7rSYooKFm
+zBwTNTH2od0aISRiDrjQVLBZ7oLfgXiDSsQI48qSIlQYSNmbdaAkbyFjNXq6Y2j
QY3HjHCyhoKs4xvc5MhsJxNtJ5w6FVfM8qri/+g5Vy1qpPmlXg0nwqAjzT5sx6Nr
RPjz6LRjpgLkQbrgzUaoLMyVPgGB2cvuNnuBxg8fVzezLTnMycqsB/4ch+0XJ7Ph
LJjVaNqRtGrhEYNIzuK2JCHRmkv5iDJIeeAG69XT9ZASvv5zvopA7U5nqT7GhFG8
romM0RxlVKdzylEYrfR9yr4k3jGJJDWOJX17hDEbD2xkkHT1rYT2fnhNnapilpGz
zXlSxnMq6UZSTd3LdxTPo0+ccT2JHCTCaXmuWuLx4ANeEnYxc9MYUUcqk3WvBhXl
NaTfYXqn7e9cI/7BnWI9F3VAJhSQheQ64KE9ZUP7DKGUOeOiNkYWtOuVsN9tnaXy
6tNGfMI0aRmfxh9FD9tNtpmlW2JKk9/THAOPgZo4MIsFdZ0QQSNgjXBmgRaqaajs
YcqfGjBzl4UrFKem2sKLKXx1QupgbTbjVaUaUpWG3E4P2ACzMMsFhwSzhWbyNL5K
NEh2c7LhQcX1jnusjyteihB8B98ImtYTRauit8NuxcLULoVA511J7O3MZKCMsB0K
ki5svmS3GpjhvsEBI8+z5AfXiuklMs/eV1ew2A4MdpQK+6/Fc2LvTo9f7uQevuuQ
7vvZjzkvvf8LEvhiK6cFxV0iBo6F7XZAZlRg2xgyrUW2NN52F27YhztUkD+j7UG0
uTrI4QOZyPyMYJbKgNte9X8xEBdi7GmKQ3+4hyVEsr+1Q2UlrjId0e0ECL7uqUdi
w/xwaFBMJA0CfbMptbno3mLBfPcktvEh2Np5/O9cNVTaefP/TOhJiuHD6OPfh0jQ
nFw5CVG51T4SRsCZZAu68Sau1q8+9PfyCDwOG5tOdl3htSe86Mv6+husXIVARuwg
WCdJZTVVELm4oU72JrbdtLm6aIdyCGcq5sE6sveGbsm/lUz2fScr0Tj4xfW9X/Px
YCnHtdixfT6YEo5K98lqQbQTmHu57uDqaCzD5FNZmXcy9nKFbyHyyxvdj9VDOdf4
DoB0TVv/HqJc03drGYemRoPVRRq15dZRYjg92yLRxJTw9ZbScrUfbntdaTxHXj6P
2aJhBzbhUxrLfu2YuQmIhncnIo4vvUHPei0vE4T5mASWk/DJfnonDZUtWgbpcNeA
t1/yQsIGVedlOR71I1tHbNgwyloiJl7Bc6CrduxpCmUaePf/Kt7NWGFC6vSEhfHK
ezP5P+zkqAAwBnhuZ2vbIs6Mx2ZqIHXBQe3OX1Jj0MYuJj7hk0EGLlglJSn/w5Ny
oLntIAjey33+oQFZd4ya3yo+M+inCPY/9mcd5/+LJj5Ckp0WeocUAT2L7414DJdk
jKcxnvDJZo5UdH15I6HuQTXjBJZYDVSLkIPEEURcAPSUiNR7PDbPJqnCm6ZEfgYO
eStTl3ev1WFmXcmDm/NvtBoelYGhwnSe+fujPkDKi+f/Z5/3mtt+M/iGt7b6JsVU
8GP9oG0N7WVWUdHQq/DoTGm5v6FFQiwu4vOfbywI6Xh9T2ItEA21Pvo0XIPUXI0J
FRDDGXRZEmmMpsFEdXUMNxZZ9654Cz4EVyJ4oZEgb+bIpuxrQMiGJ1zu7ESATKYd
0o2hajZ1OfKnOExPlJ4VYc8mmVd8jLrkNWCDjiaakh0lEOwG0S4463zYWUcEzJmg
hRFD7KmrZhR7J5QKhf68RjY0Qi+bhPLNdukMDk9f+s/dLOWlcqU2Z0LIuroCskky
T/oSzxjxDXU2e8YFBaXX3/IKR8zOS5fkMl9Iy4LflSKzXdjRMTyFLOftJ6+cevCS
aCpcHFFKH22bIGDcFySIllAm17zkYK77VW7ksftVBFwqsYwUq66H1alrINA206AQ
rmvh3PRAwgBHe6b8MD9FXaf7OlUOirHEJyvnfmH3cMizXwNjSONisHmfjhBOLaxj
qKDrX/eNaZvSVWWJYWiEYZoZTn5XW/SL3VjjWUxfWTzY9znL5/ybdhJjKGduS0Cx
bcyLUHSc8lS+ezua6Pb3SZ00OwbQmOZ+Qeg9408mNj1X1qr6itXsOQ+nToqOU5d/
w2NgzIF79+QKJEcaOhPwokaMuzfw/FaTiG5kIvKmIp2dJIm/sRfxpsYdaV7Jsh2e
N5FDtw87UMuECGQQsLuvb3WexoHxGZDL6BUkyC4IC+UuAcgtMfoL63jEViluB17T
dvrVyG34p5MQW5Y/eScLwgWS7OKcI0yQt/UPHfP4NKc8twam4uHzMnDucuQIIQai
BVfdAOYL4nrPDzyzDJXngResAN6EwBpVrWJi8eGpekQQEr+0PcETbNVwvuHuWp+H
Y/FFTO/2Ne3sakByudQA5IOh8rUdv1O91uzhzg9BDHcr2PS0U0gWeuLtIiHovRy+
XLlwkFBWrzdl3GM0A/GrhOoAmUaXBdwJ8RaKddI1t7zTE7PLKnnEClgAshOl4sbE
wACld4P4a9qPF4CKcFk/yjuJmn4xpmfQUdscWqB6twPGeZ7ezujGscmZuhhIJO4t
v4dYlq5ekrrkuhSXlNiH9AjkMraszjuTctE4z8nm1ZSWLNBuGj7DmfM3Uo8kz97A
zijGKy8zrM+fbgqzcnS/URgxy1nSJiZwA4qOjyBZFTlij5I70X9I4qzv9g9lRVgr
uiqdCcK8mrdLx7eIuZ9q3HYl5arpj9dWrtjLaifNiomqIPKcs56xUDFza++WzII5
wEpFjLd3sQyOYIvtOkwspkk0BBqDPyJHPZCoQ6VNKYaQ52KBxH1juA1USN1HXcK3
gJYmUF0lyQKHH9HYGLsP0+gWIMKgyFjWXExyz7wfmEquRmLmP1eNhMOATv1cFzcz
fGUqH3R2IEgwKOmlAi06UCL8aVJbwbJoNZ5Iyqh52wiLulnJ2xd17fGhYNs0Hjmc
+2LiqOmHSgFsbKYtXxLkqvkLEX+BH3mnynkG/HMNIQIhfcP1YtRBU9520Jnk9Rbh
cKpEVD2nHLtPSGuGWU5eBFbsM6SgOXPY+uZcUAXurbUVAlVHMAuRzeyZc0yl2bEU
ntDGdsK929t+aDPuJA994LDmu/s1d0aB5GA/IKx8ev1Yz5bI5fdKyo/Li5AbShC5
lXr4ANp2sMpqjqUEIrRc4nnPPpbph2NSZEUE7ewymBiWNyeDHSZhYVs3nJ8biP8/
Lm7rZn31f4x2U3BdMGbUSFnlgrS6+K1QG7ZHdo8Kw9bNoCStluusMchDcmwiF2P9
c6kZG++TWGLMT2QMfWF+T3jMt0tQ9csgT0N59R5hoa9c/xyHlzwOFKFUsgRaMrIk
EH3hpywN5e5jpq+GFF9FANcVhZ93CDUEWWEqcPmDrQ9eaX431QCk+JT5Ie1Ziy8M
xBz+oTpVHpv2I9GDScMHwfpKLDqCYIRvwj1hDdFdr2GVxA1XgQjk76gvCtIUIR+J
PMudqgmpfbmdwEpeMf0lRmuKR/3PHLqDW7mp2ueKewM5Mgmb4fbYSXsN9e9KfyT8
5ta406FhqXKMfRGtOnk/K5nI0AOGbWTzTfWBZ95wWlwUOe5oriqP0+T9jIEOzAZo
kFMIfES/0+6vtXKLEhx7w82cBQYPmDbaFLeMskxBeAuVeqzoaUXFLm4iGqqVTuBm
O9fB6YZGESpsDTcEhshki62gH6tmoujz9iiEj4o7Fkbet7hCE3V1bS4lu7f9uB/t
hNk/8OJwiTHFBmXNZbftCKEEiwjWOfUvXN7wObOi0y6vp3BnEdPo3vfCDwJywwd/
i6qtMovi/jpjSQrLG63o1Lax34ZXUwd9PCTynwK88A9yNx/tDkqBhKULt6FpaN67
p050W7CtFYkfYePXHSNgaYu+dKQxm6hI/rBRdsmnvgOekuYU4KeFn68+2h27ww2/
QYUSZBLsrrlH5WMNwWrvac80o2bCKuADHQfHRUXjApyQOzQFwIpWoARJOT/hNm/V
k6/rdREqwXiQx8vq0V7KM3AfcN/3zunwMiIC6DO9J7tNwneCd2weEYGBsrEcoTSW
HbNxp3pb7cfo9bcGYllQ4oDJDe/sUe6iFU265dICXg6deSYcICtimbrMUR5VqAFv
wUY/uFpyifq6JHXWlI0D2IO3mF3g8eIDJBPOnMbZNWrBakldUx9Brj9RzpKLdMv9
nbpPaKuJdQ7TKPuSBmrhh9BovWTqbRGm22zLiKIXLuz0hzD8vpg/gt2ztg+IVD3e
EDRP9fb6ZFFN1up1rcxT1k76A41116CzPxl3aSKckHlbX9pxpy+sfn81QwfYI+Am
f56E1kxhdRuoyYrlmmT4VuQNHFenNx4c0UM+bN7ftLQPwCi/iHUPhhML4I+WKJe2
7N6Wenl1wtVGwN09ouN4YfqXmwUphuBWma1Z7nVQ+2n6LToTfjADzzifXxLOQMih
zHLQGAf0++7hkFxzFj1twy7euQh0lcfgO5EZ/+fiBwk7aronzG569FM3Dk9CydV3
OO5DMePi3XtTc0sHYaHpxVukvzznVa+/0aRFMayEzqUjbIBZPAl9yG9cvN4eSoip
9pYlJ3XmUFU+w2q8HZXGB2OA4Ar4Rr5jGKOwE6dpZ4lWZq5Voj+ssgLodMVwLNtd
2eQsnk+Uqcdsj1wHTO0PqfPTBr0FfKploTuiPYLypiLCY9tfH9EHUDJv79XreJQr
/hAYisHMyGYurQZpSe6r35Y0f3IBdo9KsomAq7Kc135JYDC+ELQDCQ+fdn/3IYqK
woR443BmF6WPC7kX6ochBx5XazJjKptQzXs8/sXkEjPWyf4RTw/cTqMD96EOmRsY
EgKZULGO5DH50IVv1l3MThLDFcrNnKwkJUzLVgBGwHjua2bvL3pZ5nDhwV84jZel
dvl6fg7oZ7kYGIXvxAgq6gEqVgC2txuFzfLsO0zh3bWZfHuvR+de1L14JgcINmey
YZ2HjwPdK34bBXT2FZgWW784aWoBmeswSp30IXRwIav/guLa3hJ4+CzBepTY8DFc
m56HJ/+2uMEB6qMay1g984Cmtjd2zyJn91W1wjJqrMujjQHP3I2c0HOZKPKkLtpj
DP170O0gYQR6UuNlj7GoTl+xCxkA7cQcvct0tty9cCxbZtFOlYM4ePBrEPYUukeQ
EtjBP9hUn7gNR4++f4j63tUultiYgcaSzzhpidkL3zXg/iU1sqQtslDsOqtoiTvw
10dei3J84BacaQ84FOcHYg6twyalEqSlXkxVTayAC4FVx1hFlJbfNOfX05tx+DFE
YnJxjb0JJgEx7S70jUie0PYk8b8p6pMAjmTgFob3n8asCzUxSeqUw874ZTZq98jz
0LKBHVUWC7B1Ng2TGwJj8MTjPsf4Wi6iwTaW5g03ccVPDjlBt+6Rsey/joWrWp4b
gAUsAOIaOwr0KpLWqu9EZJluYtJx2prmSJR2pkM4qgj73xarhYDcC0DTA5jbpK3/
Rdxau3nqMeWWW1IRVBJi7VCc8a4q3O8AnEaEHeqw14Oz6i2M8YAX4QxE+/Ri8p2W
AL7FAAFw9/ZP3RugMkOHr3n9fmIQbJrCtpRLFnotHJHWqfe2z/qS5XQrNpuyQeLg
NfN2+MA7H3ClLc1uR9cGJIOphnDwRtoL47Xwe5q5N9CNSIK8751s8ODGgIZjJpGZ
qdHOTJMXW3zDuHqq8WUSyohmNeaaOuUP1xP7Wq9mGwBvK8rbfjF6Kp+KO0F8/S8q
CC5KQwAUyUinuX6puPi6MApenRHvMPIj3Fe5LPjwEKwi1RlJmohRGKyNJXVWp2GH
XmiMkg2phggabbGy8eIv339hdWdLJR17uX7gcyRdgSFFbnrz4zVaw2YC2VVTC0Es
jtXJN6d4ejgdvfrZ4tGIaLD8YYMNeU2a+XktPPRUanZFQallUQsrEbHmxvWSaiwk
z6bEAd+698NLthP8o2DFrjeYZulvJ9B5tJ6QTMncR133r1DIDIDpensPNSb/wwu+
GsyonxJLDOGEKWRuDUnwhmQXs2GHwrmHMSgSB1XLICwUJnv57d4V2Zj7tCBYr9r3
jyYiGcW5KMRL2BN0n4ySo/ii1AegBIj9qJ74WKY/uQMHfw/p8QET9NL0q6BBDw9J
5TFlFg8PP9MRKCGw3GCbW6oG9l99RxsnXC9N2hZ5Dcv7ooTc90yMirXWSqu1++bl
4OIwyqWEEp4FBdI4GgTI6EWpx1pj+bkRS1wdVmgLvRpgrdlvQ1792VN8Z8imZEfj
6KWLqKnwFYlC7/VxfBBuoKyywAMS4DT0k/O9wFBO7P4+x3i8KOWf4TG/IuozHfXm
xA28r1QbllBoo65+OLSxHlb1emIIT+rzTWa1nzglKLKQ5pkGVHmWRNcB/SX8RCSg
T4/9/h1ngO1LT4KQcudQWV8nLJW6oquLir+xJu4ygBthky5GXwXCWFzglYu5GjU2
27d20cy2PRUOAb5v0HWPbvfTj6HPAws7gpCzFrZE4XXJzHxe3/qxGX9LrF2hR6fs
t5uDHTkkW+q5ppvGAoPFlq/1XeImKJ0A6cdqQe4pkZVFNcqVPtiW3+QLoX1g0uKp
I6pKdzLJ/eGFH+mjbPfe/m5cMpdzak717qDVIQ0+t10myGZVvcResNCoMyKFcxlB
wD4YZQWb4AVz1PAInl/E7xYDL6oN5dxo8/7ZEgUTRUB5CSEANK4fS95Xqn3q7W5n
ekQpzfjWbb6PrJSrNQ+8eutzA0HgskfqSZLZRDLs3k5MDtRK22sBqs3FqZFNfWKL
zkCugL6wLyk3lnT/YMuQ28rE74ke1aGVGwldQKVbqHkuhxTgNLrdTi7CgQjBCr/g
pqROh/lWpAv+5U08uqLhi8L/Y/E/B7CXSA5XKCyGV3zhswfRo2rGol8dshbTqKjG
/ftvY4O8ucZVnFOKRTxG3z3ELrPd5uSulOwX3yB13M5BQ77LEz6MhXvHKlrq3nYr
g69oWpGjkcBqe8Ik8OWTIxTjwSC02OINj4n4FjynBdxTmv0mnON/SG6ibhSWeH1Z
NcZPz5S6v1PsoaLH89c27K24Iy1WWM2EyMTN48BUBT4R6eImstg3KMSMDGTdjMis
j9iToyPa0a7pK+B5nSIQJ37f9GQfL++fOZhl4fEHWhDxnl5qFzfNzVT1CMNbYGS0
PhErQ2tnu2/kOrtkHYjxJ3CBjWsZH03a/vzP129FRlgWaSBNC+F6cvG5cOihUfLH
9Y1TaFArkjUbTawmImvbM5t4WIXQsA+dtOQEJQTMrY6uhA8u+W2EBVq6SOLVzDx+
PNbBs+mSZXVuQ2NO4S1Nl10qS5GCeXXAcesRa0gSFkWKysuBoOYlxPFd88NGPZgN
4r7R0b/fxnX2DvqQeNBFm8+Y2jXJ5/G/VFtxCECDhEuK0m5xzT+ZDXY3Y0iENO8F
ylR9nY9ouBg81dtNmhgI4c6PvnIwY2KpEK0ImCD3eeXtJfFEkl6J4kzFaVShAWaj
H8S5GBY3vugXqCdgd0dsi+SZzcox8gamGc+Ygr/7KoxupPS2xOHeb2G2RpZaU0nz
+imk0Geh44B7z9vJ8vTNJdDT+6HL663DpDfUK0zM14iworJDFXBkTBcxxVfwA3tb
UtZI/8Ykyp0eZCfzSsfEwFjy2pb+oP2ffj5aoaB/ffWjFeYcyA7bQIRtoaBH7MT2
M0vfXMkJ1PXcUqbXHduCoRmR7Ca5uwWDjRAdr1jBOr5tYVO4aGgzer41kfDt9P78
t44ZUfgA0ZO7+P9z5jA5xG+S7n5Lk3yBbpDQ17ysEZymCVo/fbB5MVKaA7hK9HPa
1juhqjSBaQNhj8xx0NlM3ot2rOVa1P81f8S5nCT6avnq0Si2R//sH8U7eY8B3riE
7UWn7bSiM8IsbCYmZjP+BdzQf5nigzaouA1iCIHxQN4Vodtfqx+gH5SEvMOD/M5I
nqXhko5sBZYnPX7LdSPvy6vvWk5bFjogxmoBVpTWiozXPtIZUlr+fHxC9WIXAP45
UwDRQY/d0Lst91/NmyE+Z4mADryCHopJrGHJz1KmezdnJ830/T4xG4yNiqbwpey7
htZ10GINslhxuyNXlMWz7n0MMvZqKvC31vvfC/XuE8L0fO0kYa1KJqptL3xtLrO/
NSAGk1JU4ad68H7AdpsOZh0OVFAjav1P+3IG+5TwzNJa9ZeXGl/OuyllVwwx5ish
KpI3bhcqi0V9dpZQbxdh9gOgLc0kEqTt8W3WcQ/GbvjF4/MDFZWFiFpib1VV1ET9
1dNiq1Q9zMaAhWZogBV/jViOOTHl7OP+WdyP90jKI5vqyPkQKP9HxSNuQFwzNwC2
Ugb3faTL1RPF/C2XDvmNblotV8qXDRz3vUXjk5L3GqSemyyH9cZSEUHVwv3drTgf
giSNJzik2bJKq5xzjE2JbgDwVHPOZzfN0sEfR98Gmj635jXoPJS3CfXO7faNb2eC
yGTryWgjVECy96yTieNVk1FqQ2HjPIWIHVX8rCz+8oXIWN663Z+8ES8YsT5EXFra
vfRYr20fh8FQbhm3IUVORoCVA2gLHH2qhwxC3pX7U5dcxjA24WKYttfVCoO6YGLb
xdgA5DznT6C+b7v0tHODrj1X0P+rXH3mvGBxhkQfcv96UB7rwL6TUZG7UIiblH7a
sLroq6Q1E4+yIRin3uf0yVHkPcMPQrsFt2DJy/WCAHWXBdn0UM1SEFDx/qWh+ade
IXYPkLldfPron3nt0X1RSRqIJZQedApM7lkpLKVtFbPB7L1/8LjSqokWIy4YkI13
lWBqCKZoWx60j+qw9t2KBhcl3KlEi2B5S5Xe8WkswfxOFn65t1sHO0tbj56qK1p+
a2SQPHYS4ue2ql7Y3wEBJ5cFeIWIQV929snEgBG2587OX5LOQENDxHQNNWGCthR/
V3+suncPaCjCcYAaqAGwFSv5fRQAjMgSoCIXkl9S4xQotNmqkDItzn1QHsMz9Azp
ttGR+klKXK4WA57Qnq4L8Qo97JYmU+Sd+EyNJXiHifXFa9GfAb9k9m8xVgcYx6am
KUUisbkoeXDRaWJDvWdxj4k0cLy6rt7UDSJl2GAwOvfGl5QA5WieuOckR+F1SOrK
AUFDHBIimFYD+VKAIXogT9LXhOMqXpU2lzskFaLvR9YmYNQ2rRQwKxHrmgeu27q2
Gt465UILEikOgnF2hSAzWch75uLjgOI3cKr20OaanRxdbuiU9edwkc7XmQGifmdt
2GqSX48oA/tVnLm1u1CV7npWrY5p1Tca1DNGe1w7K6Orl0qiSMOYX8B4/h1JWvzd
tmd3CV3apWq33gUJDPa6gfdbpSWTtdPpSxiy7l4cipf9RyuxblGNXd4QSu4qmJOe
cuM/2Qgg2K00rCFUWfR9b1KvDHyimv4/a0xtLJi+eIzXNCqWlGtaEdn033iMK9F5
za1PAaXpiotRtITkofYClaFtCyvPsk3NhRFiDasyc1GaebH5hO6gFmH+BJhBR21T
0jU1aukyx6KmHIPnglKYwzCh6NYVUwOXDZPUyqsYZl2SjI4/5EvVoHiyy36LZtEz
UaPSnCoZ50TtI60Nyr2mxs1giHGG4y/QP8KN7UT08Jpf9nRA9YwswjiwWYfrgcyC
sGC+tV1PE4GNut6ZoZowlU3vlzqDZxwnI1MTd9nBHpIt+XiR49AyRuDlMhiGLys+
1/f5OwQbEujZSrhZ6+JkFmMMlfmIn1KmoAYPwjSodARjsl1xJdFxxwrnZ4oCYAv0
Ll3yy2v0vUp156mvHAZlAh39SKH3rAdUljV/3YLkPhaGbZZszc7PP+aaW3YiOMKR
TMUMR6taFlOikaUxNiKNmzBVkGEbSI+tiVWzPplauxTftHweZBUjVAapEApzA6K1
GsTO6N/01gRA394/KaIQzdY2CujGkr4znvkYS+EtHUvjQn9zzFSzwos43WTTmQhe
dEvxnxYLCHdnmIjKSvLNs7cQZkmusn14QWryZu+qfo90lFkWhIkdX5ZFhxNwV/gh
kN5hShySAlCY2s8NRepUltvBKJlwSMQ0Vzavisc5k1dinhbGLLjE9DqYSvYfZvmX
BMBUCN+Ot937M6Ic6cQkVbLZ87AuVZl1lxxvCrAqg3Ovatc+MVZPcShibJ23T4VR
HW0EWO53IW40YQwrQNwWWmu4NFaHVohy4reVhv3hNDFWVv4/lRuQTFSslSL/Om4d
jrPQX42cCPBpG8VHqz29iBaWVMnq7REBqolQLT4pKhKGcjr99icQMGdry7jhDyjd
L990DyJhok3N0JPmHG8wEQhK9pAyxCPh1zG/wDS9lgceK5QS0A5M5bTn2v3EhK+f
z/ze7EWa5nYxpVHHf5S78wfVt/9l8fgB3K6tbJnacUxik5cB4UgeSWdwzeieEcdW
+aLqoONFn6pB8BYuC2lIBU/ByCRSHLHA9El7f3+TrVrVhKxI8I2tHd5L6O5PAvi2
GKmU3ecuo3rkkOkoVHfOPUCC5n1y7oNRuIdPlXLgPDqtksaqo8sHn246nKF05xLW
vleVgcCRwV1FkrJkvcx3/GTvG5dnBelWwRqTGpsAITYb/WKiGQCIPrEmMMnjuIf+
Aal9R98FCo1n4ir5vlVIHyFzDJqEC4C/Y+ETlEgqM59NbHlu2EOMMrqhOiz13uGk
bYCF6QwdC28WtLKOzvz5c9RZTPU3x6qwLxy4nX3qREsQUp1XyqtshGNKuc+JgCvw
0OC72P9d5biYS3ZtooPVAOufCvBtVZ3Yn37U9DnHA0yKTeRfPmYvDPg1rpZ2TAXc
RFwbIaDNJVmNlgw2d8nZjnvL1UroMsNUhyepbhEbJCLVATHEbPFuIaDr6PFLH3YL
2/GTR/myNhtbBGPaJ3djCW7RP3OWYKucxDjgGikaccL1U5K451MTKGRj/kTY0EFN
krP1+bvYIHeI9MVEjtMB1F+0dQX/M8ROBHJeCBmI02aPvuzMmveVa5w3kKbknAc+
h/YugVs7+K7Z9idb4DPU/zUq+JWvThjVFddFG3AbRdnPrCTLXJBMO5AmejLj7fCg
r/x6bjr3eq3hU7xdW2ne8X7ujzbLwLw5EjPwzUlYxSCKdaau1qAN2Ehrj2sbwi/E
xNAW0n99BU/5i7SgENfAsI0LWZJmdQFfWHU4D11WG7QoVo3juiSnpizDscp3un5a
07FGNWcpcxAQAXgdAz1BzzzCEnLjMgo7B/nouHGKtCFu41ade9HHei7KjhahEVqC
RTkqcSTpxcSxK5Q66+B++K5WkobeJDBXXUhmEgtDzlMJRJ20geSekCK6da/PDi/L
OvMF0A1Pv8+35iCyieJek9nQwKDr9W2CTbsuNcOK/RkX1rthN/99PKYz/D5f8xmA
erZaUjMbI7rkkWdFKGGWIZfCN8da5VSeGeE6ISO2so+5tU1E4c4t7mJqerkXpSQk
tn7TljXxgWz//bKnLOztYW0NNicnQ+z2JbNUFe2y6hfGd1VSKJEp7s52vFuDtfyn
a1ghR9HkHgEXeR4gNPzQJ1JPsR1z6UZgxIFw44iMw0rDNsmxmuBA+KbuyjBAeBGi
CoMSq5hqyMgIaFCz6Qkqj7cybhIjr6Isq0MLKRyu1Y7CD0iDIPQEuSqckPR3h58j
seJPTk610cDlWSPgY7zqMvC064BJ2fILdEdCkd0cSlHoRkdnbj8feu4VbBkUYNC9
j15aGLehpAJGUlR12sY4/U4ZkympKk19DkUszBJoZL8JdZIvLlsFetgC559cndWt
1aqzZM1Gr2uSFt2dPmuAaTU3Fj0wVWoXrviNzMevH0JrKfFdGYWAyCPmEJqkjLUb
xLm2cPkPBtpa/FekqIZuUetmoBi9PD9rU8WtW103wOTZaku6Tg0XLdGfIdB9IoTG
WqdxhSlT45524JhU4FHAWExatlY/va8+QXcghG10qisQfQ4ofldK6LMIC47dGzgX
PPTlfT8lZtthPdEzyMvjhEML0G2KF0T0x/KcfG1jfP81JMGqI4nrFNCgUDaQSLPy
7R3uaQbGEFKvLk+HbF1a90qDHkrStHUvM/MnzWYMDdJKmbZDCCe7SR5yJ+0XvQuJ
mWB7snJOWBLgAPb//hhoclaVXyLlJpeKn294zB6r+uwZn0xGhINZ8aX6dr6+itzg
ggUybkV807pJ/qUR04Cg7ydJk2L7W+GAHIkTK3wXlmI+wjgFUIvNEhfrdRDBM1a6
AZMcp1FgwLyMyO05GXSXG/p/WxJjkAnqLCq7RK4c89YejEXkJt4JYaHmkdpWwjGi
s4BL6IF74QF8VwwLI+VkPBB4LF9nvQmSSmo2SfazASx2dFnoM3EWP+wUFwHYtfjv
TKE8/B6WkAZdlB51Tsx/WGp4mxduR8+Xgv2MO1Nx/+ACh+Ls0lLAdlpPoQ6I78kz
EOIt8pWdGIIzLIgbffSRCs2X0wf09umw/of+yPLEerapvbulAba112BxRmP1dTXr
JsEVeU2p3FL6tehPEiuYmBpgrK0qeyO4Wfbjb8d1Pnm5C2Z04DOC3LG0gVRoy/tR
O8qTheckt0LiPEKec06cfkn/MM3Cq39JCAUJJMb/IZ92tsd4I0YPihGmsLg/E2+Y
j4ScPNc/qwoEHBB0xVlrPg80g8CI+XPrFkHvQZ3AVi4zN00apCTL8NkVZIX3dHh+
OszmDPTV2Z0ZfKX9CxRtlzoaEaljg720TE4+A/fP5YIJULg+4NtmM1Rvnzty381Y
wwTa/X/3p5c5BrC6UlO3n0PqRBNA1nVis1+6rC2wGWLTEZQFuOEcU71kB4L8YFmw
9GJ5ejtnNQwh9fyIr1aUHl84TVgaETo/nMZCF3QxfR7HRry+Kjm3dEdfvP4nlcPt
dpMcC+u5CBv8pkOVV/RVVPeNr78bgTdPZhTJ2tcMUN+hXkUuio02CBWtOiU6xyPZ
TTU6XarFqs/B0E7C2wDq2iIFgs9nbj1dSdkAC0y/vc4VWK4BGNYPm5Fw2Er0LqrU
aUvgzogd+HfQZx7HOyRBuUHKpj2RSHx1cs1WmSKRUcc4nvhq9xaFipQQ1Bpbz3U8
CpmVd8gkF3S67D7HJlq6Asp3+z4XNVuO+x96/oqoFS5icvMUFSJXjvnm3SOu7bIW
iS7CQx7iaS1LEcaNYauY9HoBWLVPej/5YZsWWeQZ3ZU8zl0irsEcjgNQCJRTLNo5
NjGC/yIcjz45jTnGXLicobQb+Z8nyFVWOdjwdKFFAhH8931iJCZX7cZeVt+QPGNK
bQx0mz7KJok6hoNG956yJ9BGdGawOwnGfYy5V/RcJH/SacgfvEvMpqKGHOdixOtG
mSYGvUvv1R92Ox4K8ExLaRGEm0uqPS69jhSadIxD5SiB/EvpvPTKiZbZuabLxUCq
TrYvhRiuj0PLGeKsHvW53OngFcyMvpEhhKGNl1gU25xtz5p5qVhmltwJYrlqKllO
lO421Zqt70d66+TS/mgk1iDPI0IcGs8LgwT4dmPqLGvK+NIiw2iLvDiyqefANNEy
ClwJs3HuDJXD4n99g0n4lrkSuxE825lBb+B3e3Jwd9yrbuRJr9rzdxAAk7FDpD5D
WzD1JFxpZcHCzbhi+XagCFJiz1g8naTFPm+OxUkbTwDqxKt6/h8iTRR2GxU2PKd7
SQhggwbUS0gK0KFssvGnM2TkWB/QlMt0uwpMD9t0DXix4C4v7lnw02lduRfrpWO1
+pyxq6vGY9tbFEHHPOhmQa2H4WQ6RJmNeOI0+rhBDc5X/FDaTuuQa8aLzdz6tNsg
IcZZJ5NYA/iu4tIOsX/mWrhFJ8xR9mROe1hD6Ad6DfbcCti6i1GtrQJII8C6bkIB
bnzRr6/jKXejUtbKefXrN7mGLpYROYjDaxGJh0W4SATEAPwh3v+CtNDl6mCZV7mp
cFOJLFxmKLxJll5WZxg1QicAnMIVGdZG2YdYXICt4M2pL2WCATUWI+onGYZZ7P7Y
A9s0JHF5Sadl5uSu/gI9e//+8CL4ThpmXpZE6gWnb9darBcr9wKtUkmD4BqePhd2
UyBTNL4muWn4JgKrYfw2j22bJ5nTsVzr+1WE2SDvNS2KE5vXk4Ip+DlnXLRWmGXF
Q7NFUNRH7MSI5jFFe3u+4AVNAj2dM6BiXzSAVfAbS04xLEu95K0nGtEbxN1eqbeM
Te06p+DRcjQqlTql8bOf1/ntg2zCbA760eS6qg9SLDvkjejTigpma/C7y2Igfe9B
k50ZMxZE4I+zfMDK2zoCadh81FqBvib2kJ/3vrBf2Ex39xLvwSZxJt5BeHatJW3X
k5WR2GHa86kD4fGJrB20zZ7Ca01gCOBFhCHPMZOc5hyNMvg6we0G2jqrvKUbPogF
l4bmkApkE14ecD/qoUbDHjKte5GuLDvE7knJC+Ujfckn+Sneg9SVIYwXR64uMbVy
8isI2DAA8ko/TljwBJbarQGGVBbeaNf5sZfiSUvGH2XW7ut/28cK43Rk3sHfO35S
o5hHQ8Do49OhiOryZ7/3bJAEfeD9+ARMO8i80tCb9EynXTY4tCsSlZPpPDvq0YHY
7dgBrvjmvD5g0M8yz8c41BLYaqDdSeUwCeywaffXWg8hslNm0FTglluta0YGMLq3
Rf/AyvIg5+GSmnf2uHtjEIETjdTB0myyh8U2nvslGEsDADT2Qz/xNv+QsLNMV+id
Y1LBbI8bVjuGN5msIunuPH4y3A6Q+6LQqFB0kXVn/4qtd7EGRCzbggV7Sm74osnK
S7JNP9QKbkDitnQJAws1W3d69eOil+hkJ3cX+5I0SwCydViuKmZfnKO+F0eFOXDr
tYy9jm30OAvHMPrni1wCGwcl2V2k3ulrEtG0lNA+++YneEZ+Tmg2LtWmRV4ExDpH
qBTYql4C088q8LsS7x5uQtsr3VaZO6SERaorT1lXbY/vvI/+DP1uc5u6B1gpFMjn
6xQCYlbD9HIm94Vn6qjWQwsPhBXvYbKSVAdAzgNSIsY2eAvATyz+Ningi3OJuzf2
qzuNJuXk0kKVoTdh13KFs/lJ0j3qUWvBQEz+6b58XhMtFtB8yloEyYeE0zGJBrbj
P1s8BliduprhGhxWecKE9sYmGuYuiWF5mHm1x6+VXSnmftQId0w5TyhBHb+R9M3v
P92mR6JFfXEi1kUX1pf80bjuhlJRYpld+nS1/DEsvIpElkjUTHzfr5i0eg90xZtk
wD8q8uSLepfq9AtcYTu5D5o91CS33fvjjXuKqajW7ggApKXHwHZPE9XHlIenvzPk
YAy4W/f8lGEpZtEku2jMXPyOfSx8r92FouU+dlh4VixPFKMXJqLFRE8Z42AiEMZ9
wpSHxT2KLdg6t4hltpjhYq3rokOgDy/oxvFP3wiIQflfP5MVj8kcDOLl/C22yRZI
ZbnPP/KP4n219ITUkHl+1RrzDUD9K9X8kNmIBV+4pESRLO9YU4HqH+3dlh9mo2Bv
rbbga9kdmbQHp7TsZrTfbXyuYpR4OeObcPx4BlLl3dHtATsdEKCHrZ5KzIvqLg9i
WapS8EVzB2U1rXnUJbvB9hUjQKQ1fA/ZxLu9bN6hT67agstOFPSsIa7dagUsi1wv
5rGUS4gxb0roF6gGKQW+EpqTNfoKpO8QLkuqXZbJHBVclojWjgg1WCk4WP2Ir5DM
m866+7JsPbh+4KDoGWrcR8RxIUd+RNAUnjiTgb3uR3BBXgnJuhMKYNX/zzKWa+/k
Nnqe7i+2TOVeYKkkojDMx4/p5gsWwxzHlZpioSwSx4rpf5n8ET7mgB2NQfMvDgbO
vDNqf4CLzdgiLzPJC1fRwpWLWwrA9c0phpawpxt5M+ZNH6zhJ3kPn/b3KqhPLrvx
Yq/4agCJQxDif3/tRgc+NCN9D+11OCL2YCvCHOw+h56rJWLrVFpRTQJkWB/IDiQf
N274x97DDUaMdf++q7j/g/GCE+VjT92HSXdk/FngSCjPvV7xfLuhxXTMZRE9gzMO
RxJTaalNw0+GcmaMKDwjmi9qRTuflF2RlepN6x5GweXIsNeq8Fu+ALdBsdUZ3IqJ
bh5k14jWREjGkDJOlPVd29zrRDfQvi+gJxrdJW+jI8tbbWDfpMmTrbqqdkp1gOtW
8mAr5Hr4F0mzsvzUhG65uw0HvT9hPDuoArxsTD0oJBeJ93cKvvrXMPs+nSGx5ygB
xF8PGFUE6Tc+Ec3zC4+HKKflQaKoEUXLISTjjZUa61mL64Qbrp+YAOs/+1mxnwgj
m6xVfjl0hoyynP1inuEXhc2vwHnD/5kFqFJweWm08z4/ZIWqxLAzQaFFDt0uk1yD
oq9amPGsHznWkyZ+cebJuy/OV4Yns+6lNv/+LmOAOg+xyWsnqUKRn+NE0jd2x0+U
Jvgoq8YdKEDuxR4WO82poGH5NN3Mg8OMXaQiwVXNj5aVzx+SMrmzHxfIXm/U4r+f
K0P/AR1kTN0cAng/qeOU4TiPmcIqwN5dy01KKIotmQXsNd+mUwjp9EA969wqKW8e
T+OwcRp35iFhszuePwlHAKhhaKxO01wXNs3j9WvyafnN+0sgyma2pgst6/r/MJEp
IhPeYwNosyOJzBcHQoQC/hQYdW3IkE34BU9lODY+SlmXsYr0oe6Pn9uwj/vBEphf
jd6R1xZwI/EbjjUS/cNJNgBECf5+NthR17kzna6bzBqoDbM0hoh2e82oG48i26Ti
1pFdTDYO/4xAcaLfiTzalelUMSYgYmsUHbGp34Y2XCPvWZcHoSIdQD3rYUbeZ4Eo
MyP+UmmYvJz1lcrhmCNUwZ0LnnPIjqTIpcE+Ds12XIKTR4XCoxYyyuKIRnuFRIJz
x0tYXVVTpJeNKfj8nbbGwHm+vf+p74VXSjNtJDgmF3+RvhPLwYdtjn2ZQMMO7DHD
g0wT01e1avzBzob6OWi1Vibb4ki+OZHOCwvSYN35JXHEUu2EIApVtSstBVxczHPB
c/AlN6lLInF+cSCtg6ehI/TiZNK6St4rRdKwyIzReeo=
`pragma protect end_protected
