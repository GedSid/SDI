// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:36 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EP1JZ3pmcKyJsYt/mf4xfH+Z/rJQUZuj7YcFnjMKMQEl8M2n4h1l1Vc6PJoIrHSD
4TOIs9t1akbtOe9lSCqk6vC+LJ2kYH6WEBFeryAJ839jCymgqdypV2zrp6bxzFtA
Xxvllhvt/IjSSAo2aFqVOVC2sd4oKMmn8CL38fBtNKI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 104704)
zuYAA0fvvTMS/U1GKf8TnXqPqwtp0HzHRNrgI1af6ys+hL9bOoX4SbrFllbMPAq9
CGaNCaejJqyF9MBqzH5bz+vhy/HkctwHJ2HBlmH6pP4u2YOTA5yxelwybnO+1jbu
cZwXgsjyWor5K6Sz8dzEVA470SCT9i5jCXn1sSYHBMphf9I3E66JPj9lWZGZd7LR
d60YG/txrm6gqaOVqcGB9g21jpl4eP0JtDMctYjic70ZqIg/j8v+F7Y5iObrDyLj
2QIuIisCR0erDBgvPjAFT4rAhrMwrBfGy9JdYlh5lKELTuF65MsUKmGBqqrm1MJC
CTZMxQn0ZINVlk9hpN0Txvdh7vny1sd2LXLnaFHjw8z1Hv3cTX5eNhLW+Jws26mU
AmJa8fuGpp7dCbRY+LuHgaPTCvUxkqKy3MN04DNvKEdYBdViFdf6nLmRZbHha3X3
1lpXAhqo5XmFqs+Vfa43mHngksCryzABQc/L9lPTMX1nIhSm+wdilEMNF34zmZg5
lViGHVuu5M0tgPFmTOs+DH80hP0LLmJ5EIXGnBbHbGg3nDSKX47Xdew+RCe5VoDg
cCMmldiKok+TwdkjLWpXFlTWHH/9ELBu4MXp9oJ3XQusmdjfSj+JUPY++OlYnbLm
kHmhXCwByUHJhGAso8c3EbM9p7an+viqYPCGcpSqzk9dGrZY2LASIB6VXHecH9ab
vOHTDrGhXRUf9RRsr3qsrrfJCSDo+hXntBkf28afDsWEmcmAax7AfqEAHeR46wM+
QdIRCW2E5OgfcCFpg60sZIHf8tN6KweaxZ/1arRSRSzQrmVCThVcGQpXa2Evf2OY
1yh58W9LpbV+AGo9H2v4bav1wfYiJIMCkcL8yNRI+vIPrCkG3HYwMdQlhKOuqN1u
0nlK9TylG0Gcd+r6eRMfmHVUirsohPhLUcBxqKOJbh1siF8vHl3WhGqTamS0/xHX
muXrUbaNhJZe0r8mUEaV3vH5jTQ+OuQBAOAPd4HtsiqGj3enGoDkIerfgpIoDZmJ
hBuTI/5WmTQIeHSa8F6OerpH+bRpH4FrQcJypVLBh0we253Lvxg6ukrPd4CIgPuz
fhqrADa/cMDhpb6gsMYeiyeiI7IqUpUwjxuTYiZrCb249FjH5nb+GHDu7a32b4yb
9QW7ZFvfCoV7VdDxktI/20+9kS3nmxDok3ViXkBLg7qU6FHjYALcsavH9YNdlYUe
dHQiYsCPCEarAhr8DQhI+noNZbH0UUKOEYSWzcu3bRLnf78ulqY5CGi1Zu5QZh9d
q8K4R+nu5Gj6hDDpj+3A5F3ODOv97O5efZpQvY2qrqsb+Qn8yuSwqrvbuR6SbYpe
hW/m9f05QnoSBfPaoz+0BurFxu66TEegv4lsS5xcD6iD9f7sMV+WbIKAMFuQNmfT
RCUPRTK1hFgR3GdXfG5QfIyGr2x8QebhihTyqZdvjRxqhCyXgnaFqMNJTL+7X0lG
33g4UDOOjXPZ/ablNKk4zVEtG3TINQsHFw3Bltfk1BXSnA2A6HRc/UqSUIhuKsV0
b5UTH5jZfvN7WMKA7T3ZJ/qdHrRULeSVJM3wDhmvV6NuYgv0wu+WTF6+eIR1qhTG
JAV+Wxo3lpv2stORAPrYzv7TRUJlya1aVeymFT4Q7Im7gLraYE/E+J1JyTCGLiIY
aTbpbwDEGOKq0xNSYenCXQXUjxNcJFOCStyr/tpXiH13cfCfGBMTvUYmlbbHUVW0
vVwdHCBG4dmmPKDQyIJX/hZTWkQZH7q4UBF8fZgTRhD3UCyiB0/9p78lk9Oe7XBy
Dih5JXCsrwshVG8ecY0sL5yLz0HUaG70A/uFfZUl7tN1bIVCO/iop1imxjmJSrnu
F8Ae7KZn8yrb8puntU9h7WiM7uIBm5wjWff6+dqjeBTb+LxCyo2R2Xk6mC48UnbP
HCiTUaoKcsaNaJv7G2UszwOvfhIRHNItjwiEMbEh1vd/EHglhsnOIIGfaMyj0qiX
xsX1nlD6x86y8hcRHyZz18ubtIemyoFCYMeBtw0wKzE1r+BUwU9f1Yl7VeTKuu2r
Bjpx2LuI/bsgD4Gkngyn0HpP8Thf/vYVwevbBZLGF8epLTGFxn+nHlsLGDX2BxvC
fgWvG9z387e6S+nkczxWslKYNKCzo1srByY5rgfDia4N5RaNfsAxOrZLV5NEN+ni
0/fadyUfeqCQ6mF/gG8OcFNa1CGzPA+492V0CfMnXuc36vsj15n/GFeaUI98draV
OVm6M4MSJ042v9VoNS9ZSqJX6LJtmknsT9rgo0c73NQe/bpPoFZ8F6UhNTvk3zrO
d1eGFUpR464xhKmWhcmXrWOKI8p4974bl9fFCnPz6kaLpLlj5BxP6JC3ZbbBhPb2
9lnWAQ3NAEhTO/FMHT3rSf1QnTt7ietQu7NAQ1NQfnXnS0xHt+ggBuGw1Md3abVW
6BM5vpWSCZEJ63qnqYzGCdT8oSRWKR45iHa0hkzY4U1pEGpOF8FQukJdr2x5NBiy
J3uIQOcMy++lcAnEqMRyR+GeYzvsMevyjBt5qYw184b9MFen3qfFOgnD3yfR2xfG
m6UDJwh0QIIYvImwSJ8D90BS+T8c12JJCIlo5KG4utON/y+wxioNqlXrwkJIvkH7
s/CeKpPRxvTmvnOKvl5kQya6KUl5Y9WImmdGRFuk8rwyiDKdlwexYCpdfXNDC4zi
kD65DIsiMfm6iHfyjLBiBsnGqm6a9l0rsgqnpvoJOUHPYtuLyOlzcDeD7T924EFM
mKkl2hi01tqhzsaakbcF1LqiUlW3CXY6RBSFIMPwxk/H9zbd/A7jMeTXsE0rs3J9
3lyAvu5BB6LBno1Tc36adSfIjpJW+UHWASxEHsP3uYc3+pfQCD5WM52xRrfjIN24
PpbK+EeBmJXzNlYBy4py0iEn2jgb8UhH/2ip5+fB+uQdYw+zd0Up3dqo3eusD+n8
rw2OgyI3Yuarv90kWii41qeV0JI7GPagaXRecNVTc7Zu/BSbz51q0e4TAno1iZVi
/YiLuyitQlK9Of10dXQDGobZ+E5/DxEpXspToa11lwGh1tnqjqKrK0ff9CQivNOL
OtJn0BKS8dBRZ45BPscqJ0gPiplZj4sff2a8ZyHg0c6o85hHEc/Vdb2epvPHiGmx
Uuw5xWe4Gdtsk6R9qLPjriewQt37RZuootdLu9oBDISWv4T7MueVyA3bnsOLnEz3
fgcSWIw7rpM18DxC/pgTOPO0D0zO0Mq3TS8rDL6AUcLnUaZTnBsqTfjIF07SBERj
qD45e32i0Qt8u0NH8zp4YiJis92h/04dGdLAJvgYYG8XTaTGZMrOXbPI+RlbPhXi
JCvJr7ZQnaMqy4Whk7hDvP866hCUaFu/39e3vwcOfHfCy9uVHL24pFs33v8KNUwJ
wEKMvii3ps4N2A6Jakwt/R7JC7kAzbaczgOkgJQ9saLox/l3aFJC0Qqbo4ggnpBx
VQUoJqJeEWG7N6b2OciVZJ7KLhTo8dYWEi/t61QUNbwmJptGJoO8Mc+PBolpkpeL
Rc7GJDa8JvyBtA5oi7/EaDc/YdrfTb05KLYaBeg92SY6heE9zjDObwZFY4bvYghQ
WOqhBqksqBRunfAvhT67hgc0Iq2kNLsZxakUTU0XXwGIHZA8Pdg8XHkp6iyCjKaJ
1cl+dqpY00TCc8OwFnHzSpOap2wZSLdVZhRES5uggam+lNZ9D6SRKJ/DZV3UvvY+
F0f8A8AWrK1e+lTEHhWwEOudI0xDCwdwjFYWrwpa7zkqqGBGgQpodm5RBY3HFJnQ
ElZsUHvBBC95JyNMl/tS+keHY86syr3A6fP6oM2cX6zOOVPkZHPs4/ErNCc9bvxq
xYbfIWqEk7RoG3tSa5/2I5mpX4fGY6HFf9LBTNxPmpflgD4RxL/KYa7Uym/ytqUL
tAH2e1smFancqUItv+nVe8mSPnfAgpFcnBcT6zlmSuSt62TtMimbM7rtR2O5ayaQ
E6FXygDoVY/+6n0bucEOWVj+nGHE63NVHYF6DhsDcQuIE+WNAfgLnwmQ4baR0Ey0
015zxV+ASjGRhEuCTOmDponGmdrbHWrjZjpVH9bgd3Hd/XIXC4x4VieURZPfmUhg
iJkQ5iTnEtUkolPopnvTtAwKTrMDlN13EW1S2q4YR7h42u6YvMkVefinukqB6tdc
Hdm/xCBUcWvcGxjZ1yGj1GpTNbGslH8TuM64aZWBhHwv8ElKxtzT0KfZfq5D4u1S
oIJY5FWXVYIcyTHqYHGBxcHbS8Xu7WV0Yahw06HrYgHEbFx4/40GYTrqMKiCb+l2
FkrRCjn6exyoK7xqPgHleMrjb7aqoxxSJGy3DViZKmSGavWc8QhQFt8QtrtWaZIg
oOCmLPL2qWP2mBB3Qtzvl4Qrz70YvQJcaqVypDk6ENiSOV4D2YYMVQYBsT2PA2NR
x1MSfuqXS8fKpDBTu0/az8cIUgLsesdOAO3Y644m5pwnzwYQh/U7ILfQmmfZgU6K
kYUq4Mxpzr7adcVOFMh6czYaySpVlEN036aIqoW8XqnEDpttLN39abFPbXR/2X+A
3EGtxKSz+E9V650/d0fpMDENGrbxBUKeIjtpFWR8AwTOGfoVltpb1OUg2DESEEky
sZGBopfRSxe3ZVnlzaPiq95F7JobvAS7S9HV5OaLCuB5EhdRrDvOCsWvPLNXjUab
JzvakgGTFqIzwBUsUcahqmzPP7ogqMbRSUMJHVETfJ9ReG2PYHAprzph16nYHdpn
tLwA7b6D94gc8WoXWKp9fOspJ1R6wXCf9npRAYVM4/RLRfg31whIdebyGTo39Q7Z
UU8oEweKxRcAbytXPPGGdBxow6BINIo4oQptjn2L9ZEdmRvHCnRKAR7GfD3FcjLa
FrNsUnkJXkEvlotchptRwy0OiulArlY07bZ90EEi5RlFs/fJh+V/rtUZ4p2tj1PR
0y5pmn4WnuMt+pgUpXbrLuBqEPEiq9LjysvazAv8Az7lOuyC9ZWbJu+sA7OHjKze
Y3rs/pV0A8OaNHlMBczn6tGi7fw/BtxBkweSjX9GfH8CGUelJ8IihIwEzjTrWKqZ
faBIGvE0V4S1Kwqb2HFix842DIFG6Lz2wJArbJWae5wjOh3eptuZkz+MqK82aR7U
U6Zp5S0+p1JKL/SoZCdS8SKL9+xtmVaVA6mlloweOe8Zo50unGVn8VOCqv8HU6rv
OOxDagGjkvJJMR5UAWFjwM5vmOAjrq8Q5qsiTrVBWbojtjpysC8sqsFPOd7mkfvm
EDa3wtNPKKrofLjJWM3wt9HUoKnDld0uL/yCDDLTFQN756y8HoNTnxkS45OMg5tl
T8uzkxTVMVDuuTLnqZBjpCjsRNPV6pErDszVo6bYlwTbkwvedg0Q6EFdRts2Zsxl
2+BlEaxxznyYO0H1iw4pN3s5Tc7i3RjPgY/GxN6p26e4qejnU/CsL9LsEBnMFmRe
IiWqZih0FmyB/PHzkLwqG1daFA3X8s0Tzp/VT8Oi4+POfzhkWHHFYttWYQRCFEs1
gEbM8+l18T4nMywMr04Lqth56RGiIJgb8OtkVzr/frbwRixc2mwPwwLi+dci4590
UIOZaDbJW8ehcHH4sqQIz/0G4sdq2jJ8V42TUPuScqqb6K/KeMCRNeI65sW3VwF2
Zosm1q6X5cvH23BHtQNZ78Uf0KUSqIZr46yn9069CnDJe1VlDps0YwvU35l0mADf
EyJrfEhLG4DtXlS+EfW601qH2IWXjAjoDOyWkRHxKKTfAeQWhIbCsf3hTUWu9Qne
WVWQwgWU5TU1/hKXMvENiiNcAU0jX7Zai/OYFtS+7K+0mS/WSEoX2t3V6KRn0oIu
UtfflFuOuOY3abux5jJu3ibp6/8TGz4t21vZlSdzgV9gcD3BLyBIa6JcxbbvDVSV
xNyFB4Xss7ZpmXd/KU2Thj5ADZ6YOAC6EqgfZ6Idmm68Tp/vmlpZKXM38sOV28Z1
jb8QFQySYNoiB6CDM3OAL4wH+3u/17STzM61aCghASkKo4pDlOvLDX0ARbKyily4
nfOHyQw2+A4TKwnmWDYaWiBPXbFX7hdctt61vbccuJknhk0ZAsyFN93EyV8Z+fvt
GU0zxdO18K120gOnxmSok+yYyJA/J8A6wjgNFnJF6kVyYh0LzaGHWAgIlwiI1KgC
yB7Nti5Pq7oJWKYwUb500UyDNQvd9YpBcjFYwK7ajLQNdb7XIoaJoAFxfd6dHzCa
/aceYXRQyxtb58IdzDmSBCDhLMN85YcxFF4D7Kg7tiHBzH75as43FAYhO0ySRpVQ
Pwmdt1ptO/Fk94ebcWmq21JDKQy+8nDQRcIcfssuaYtjybxYYImYc/B61jY4WZze
Jh35uzu10SgVwAY/aHoREDwKGIgS7D4oOBkiWQuIV63QsnTxeGQyhMVMGroAU4nw
dgSfz7thtCTIXqsuNCvcWxZwBgEZr08LL/mGZApgrcEZo042WtpeBquJwyi9IpHl
/soEL+M1uw3AYqWm+BMjutHNOZ+oGcNTUHoUSwZJ0iaVvBQ62jiBByXLRMIWTnCk
WTvWXZuDH3jiW9YQEJrsqAEu3h2TMcqSj+sAcwcJjdukTPwQyMpg6kDzvCgZIR8f
ovD7kb3DNIZS/cnvnfGw3ZWQfKMSPZifkTCjdTOQKHhRUwEZm+OoLsBvrOm3ux2U
sEt4Q4sZpj49VV/H9K6IjfjIBSXog/6dxcrC22gtsWc1xvAYcmsE0FlYSlOvqIAq
Cj/dMMLgGT87gk5bofR2o9TrknmLrIK5lcls/EIWd1TNvr/do8Ci/UhgJDyAh4EC
o7ceOiUxVUJK2C1TXSqanH31hFXV9SzA1DTumuNGL0Gx4OpykUIQEhVGXvcSRnPr
6ecPgmYhO2Ba9iwby/6q0Fy8RhIw8SHfRRM3MxIdWqVmLtZd/H66W7TljmVjrzsN
NyE2EZX6TOydBBlzNK46qNpKhnAe45TstvGHaO96sZhlYfELFp7gCYJvfBYGTuIT
dI17pCIJbJF5IoD77pmL3C9CJ0bIALJsY4SiO3/sLvCnAWXEN52tvW5IDyZnrCCX
2l+ya2MzF+WhKivVS1Zmrgf7Tjd+KKkWqfpbvdwi4egabcJqMvzPHy4EpRGteaSQ
HNp2pMBjdn1L4JQoPsuDJi3ow+MO1kbSWyy1AL6g/6qQUctpA+u8ZPxfPOsoR1Qv
/wDlfnjAWEz8toGE/GEt8MejKpHdPsMMpMdwkPNQwD/wUoNFuMzF/xrt71D7kpyS
JAI7Ib78CXg2u0j5mPkp8tE9m44YQAAlrBIXjihPln6jD+5fsIsQ7J1Pf4nskVWQ
9HDGi8SkM7ufdeuAAzOWaSh8rG6A+mXJ2j3jPwH++QG0N28plhszcY9go8hhKmYL
6tMwiYYHZKYa0zl8SdocfPJqpfBk5fjtTol4K1dC8jEtmUbwHBwsxF4pouLE+KFT
VEyMGfQijJIkVF+K9cFKa6YFz/8U9YxGjtxSGFtfB45zhxcfDDQwtYFYPvXAhI+1
KOXmWNCUJcJh3Xeg/sUYUnWheueDLU+Q+EhUk+Cpb+qugdbP4Pwji2r6XPWbJMv6
slNx4IZeUyGKnDkyX/53+DoEFOEjP9OjfJcbbslp3TJZWUK3jdP21XbySALoryrg
ABQvKbV68jTwnCB/GtoINK9EO7O+HtyXeT1EYF2NxlhfldeTMovWFl0lawbzuov1
uRFG41vzZ/DQ5whkuQ25dx7Z6SZrBBgm33iad7Y3HWLmAJFsOjSnx2yucEaGgleC
te38/fo1BQw/g4+Q1zTVyA/bESbISahuzKAORWIkAqE2NGkupqoMu+FZjl+FZHeY
NKR99fQBXiNyqq/wFJDLmCjvvd9ED52e6z30AQoi+PPo69Z819Hdq0VQ9C1fV1AF
cqFB28WNtHBzAS56W3MhG5OcKAXPMvlUumWOuG4sv8W9WYBdtVn4SsRKzttWmmQf
teK+BwVm4zNmAPKyk6L+D46YtUqTkQqmIrolyjqWMo6+iVmCzhRPFWMC7B8PLOGv
hdcMQ1ohDJqjMg+bjWVR0jpIB/eAci1lBWMaCXwcfy4ysmFPAYH6R3FrJtWcoI1W
OBJD9c9rmLAJOQagGelCLA8m7Zl+6AilNS9B7J3PeyfgfPCu3v6GQwZNGHJz4H55
gEB8S1yChgIkAp9V5CiyQFFLSs5xjJ76iUGgLWImV+Le17rY0vuFiHpA9rHxQ99v
wOlzYx5BXJK7Aw5OaUrl/iLfuGpNvAfCGIZHhofHbvwc+wCDD+uPf0XgD7fbQOCA
QdKruRGRrN+fW7fSB1/UZCvGcpLLicYprHY6D+joS1+kHhHqRPXFN0WyHtkA8xXM
AfRFgWKyUR7/32Y8AMfct3kfqJqpTuBGlagO8eLlDRS6AU/oiYi70USOfbU+NxdM
ZU/eRkpFp8AC34zVhY2s8cOwi33dL1hLjahaudjzXx18bzZm1ESenNPQHhpJXi2q
6x0Mu1nalf/bgMCIso/qBhH19BAoc4/faUn/p40/qRwM+VnDfeQmithCv5k6Z5eO
Q3g6UZ0kQlRs5+gi1HW8wDDDwz1jTTuGWxxIWSldPOA9RLyj7ssfENf3OIxw8eTN
iAnTfhsg4XQIS5GPjl+eZfUesqBIDZVGuVrQab11ZMMoYeKwbtigQsBpJZlitHCc
Yt9w/Hn82WddTe9UFq88N1wVpAB1FIziYyrIVe+2+JVv/Y8W17Kn9XglWaYM5LiM
udpMWnEwICk4pthJYfZTlmHg4bnUctk06a/nd7Mo4rURANVk/3nDJPomVQ9E8hfo
5w3+cBlusS2OMXOKG7C8UbuL/MEknaKI3ntBbPcMRR7ofH6QErKoeYcQYmVHHZD3
sop32+9mBfTMder2R2NVQdjSNGVs4BLKckIPtGEVALaV4yrzuI6UTcEXGWyg18pH
KWxW2T2VtYWm8lWAF3xIu5G/Y48Ywx56M5L7x31jINcSShSUWPdzf4EomyJp8osk
HI9PmnUz0iZr0fGKW3Qc+KvdlZjD5BE9gfIWTHraGV33dBlhpBdSabnDJug3cRWi
kpFr7utnXjV0Ju75fOlaoRrovp8oGTVABcOlZGBiqA0kbgJnTvbt5cNdBMufARbk
M4GSyCJF7x5Tg/tnD2+UCTx0hOddtXnSbdobIW3dCmT4cVeqWNjUrKOIkREafMBX
lDHNHYFoKEgTzSAYwmnFkBzuOQk4StL7TQlGB5LnqA8UiJwuFHWKA1bR3XuZm+YH
gsvfHsKFc6CDmBrCC4m6TZAa9tonedMbHdAmWlDqK/SbdXqasq0AYxyxQ25pmlEL
RUDSAEY2sbFfgO0RVUX7GDJ2rmV/r1NZkZuykNrsHEpJzeYZzCyXic6qTbdYGQ9/
LPvsZaQYY4GTRzIrMXoNcUwUNVny6Wq6r/879fvl6veUypiJGfSmfzVIorYZ5eQa
qQkYBEAeqvnCAfRKSDqt48/2Gf1kZrrV2hbWmmgs2Hha41od+aN3WOxb7fFcVopF
A2SWcOy5YMm6pJ5lHnmDFWIJX1I8kH851+3ims3fjGH58DmWn2kn7sq1IHqVajZp
bbHYLMFT4v8ccrxLy5FsHiNy7/mqdXX3O8efTmJnV/+6nATNVjxcv7IgRf8flyne
UiN1kvaI45e8VuwwVQmVX+wG0ASmYgyBjPERm6R3WOQsJKf8RisZeOsL1/Fw3HfE
yQyYpU1oY4RUJzFltIu5JnZeb7p8xwlyRgxU502Om1z7/44RbdF2AL6ph2sb0A08
gJL4uY/mFBI03P1qbtYmfSAQkIOmSUjgNMr7McP4IMtZMY4XblJfsRKjRGwVJ5am
w9lIjtuJRrLl8lc3/7wjoS5L9LeuKF61r9F3gryUqtxpgoLpNSyncuGzHl3t86M4
pp+66N6iktsUfpUI4kH3xZwlmvWobvlnIuvX0TQpluX4dOJEtRKOJ0LhfcZPer9i
1lcH8euIXd3/yxhk/zouhOksSVmB8tOZ4QylkWrE3jLi6ZhvmBB1r5PXvBt1EYr4
/IemCM5hHzkVVgx9DdkzSpOzgEnbl9L8g5o8KyBOY5emWaSJNTUS8DgdCeAU5bKg
NcwueFKY6gW+unMGfN8Rj9f8rhndU6mvijJObXCOZmEGkaQNiB4ju4ViJXrGJUZv
i6lwrfumV0et1KaVH7is5iEI0eBwB2k1rDlC5/5oyYtwM03HTxH2OgoG61Cy9UAs
q6ZaOgyirmFlNeWAnH2FXPtpX/8Nbr1QEROXC1SXaRWDxGU28qIVwPrFt7+1MRfG
XrAMYW55iduJjYzj2KfNGiIbnL7wmcjhvr+AjWQyT+uVsDLLFjsyVHFYLQ16M3ES
S9p149Ack5RumT8KnilPM2KGG8ihE9R0U3ZGxMJqN8Hk1YkNi0h3MU4SGo4ir1At
BpFkM5sMKG92etp7PFoCmRDWSqqjczNrqgI4WKeJaXm5/e5jwpuxVTUQ9GTwyrfz
Bbm1O4WYCYYPfthC1Ck7hsFX3RMwacETzgGCVKPwo5zWJnHc3ojn5OSDQiaHOoBj
QDkNN118P0Upfkwnk4t9swRtQ4jLdZvdCVRa8FEYaN3fzQ3loBpqyjc9wNNEdc4a
4Ylh6XlAD4DoWfnCt7ejA5IBCBxteFALzfT2qkpdEJEDiiFLYSNkLilS8L8jYSYa
9aPuy9bySSVIQCkG6vTcBQvQOB7KJPEXGPtz6YIMB0CcRnu11PDPQieS+G7rHy7H
5VRmQCyy/ikK5cmGISrBehrDbxW9xiU8TQ3BFYUgVKsoHNJjNNOKzWVWu7x9jCta
Jnj1kuT7fwOVU2HY3OhjeXRghzs8eOOEKRjegP7xIvm3n97btDi0Jl5XMO6gOPpd
P93zycYzqLa2fCu9Y0ycz2xp/5SiZ8Vg57x5C/RyYkwxyjkS003lRQwpTfjeHBub
evVcGE5Hx/HTN0rwRg02Vm2UH0n51euNhWjG2CMEo7dcTBpWIWWI2tbmAVL28ecr
GF2lvWnGKwkbCtnEdpVofkZMo0ZuCzUimEINcKUnoOylaK8Zqz+3mmOuSeVjLPUS
0RfdRv9OUgh5xtDlqW/oMJO5NmFSUnmKSFwF5m0IViNDAMwteeIgJ602th/qkWab
lVvCEsUmeM2Pw4wuhNOBEGNdDYqvlBoNnElB+qtOEorGLm0mF6hPbomMHRfG6T6A
q2bgm7uny4STPpMq3uOvzHIDWVd2B8TrANmMJ2/LGsqcoRZCE8c4TgDJwEDGCpeh
MYtLgTzhjk2qttIGFDxkZZ0tLRz2TAaqhb3SmVvnbiOJsVgWHoF4uZpWsSh/weRy
Q9TKugAFDB2QTKRVNyLxdte38twA35Jwem/0VAjtpzjBjW4u8yKq3ygn1myFINFo
pwmdbsWO7ZJ0AV/efPfj4DeVk3/ZhOb3MBTMrII6N8gZ//9ssqFfuA8kQzqaq6wc
V5HSwxBQ4hY1wjnq5Icibq1oQrEGjokmLy3oD0e0l0W3SJgiZK5c+HL77fOZsMxd
6Q1fU0bi6YRDj6xijBMAh+toCQd45C5Br3BDR+U0/anh6eyHSD6QrHLFeXzCWc+w
HEwq6+WMNdYj0JcdXjC3c8j4Xqwdr6Md3muY5rVCx3j6tmoO4UxzHliNW2rfkIgB
6jwTbU5DwRP3TRZWD/ONXQqYOz1J5PqJXxkMsghgB5y8oq79iDVs4k/9j6cBqw+Z
3Y8k4NfHLco3O+D/9qP7Ymb9FT6P2nPoM5knvEOwTgc1k2QEx+frwOyC3c+Mkuou
X2DhcT0CI44vQETITtxsNZXa+KlVnKyI64E5734k4OhN+H2LOXGPiBH1DGC5NerF
mTQWHeqOPN8qN4zoWr6jPh2Eza5TtoPmuWTh+9dhJL9WXazfnPxBt6XL7iwjJUVP
Ptxrl2SLMiBKM8dmKwIBTkEzhju8bp13lgtxOGf/XvrSJBI2FwpjVD1duSm/0hXK
o4a0tF7zAdoJQLm+oS9mcdV9Ihn6+SKyESYmyDbp+pjoh5gPXLSDzeLKsItGcRjZ
E2rCHGtZz307xm+NwfiqRRsbujdR919UyyRMQyYBTFQeWWK0M9nnUdv6BdmrMZ+S
9Lr0GOp0bEAEXxSibOJEjMvpwYq+TZNN3m4M2ZW6J45O3TKa+ed36W6xwBjsdM5m
OYFNTSHNevilq8oh0iphRqcPY1jO/VEr7Yu+NRv8UmROINPvhALhSmueSGe5kfce
w4o1d+9GwTopdCkmnlW9aojEm6m0DpHnXaNFFMYUBT8ukCX9eA3BWd8nETkbD+3k
lKC0olyfySDKpw7NnrglPhWNMovmRhryqf6ZYCBGqMaTv7LfOODWhMoWM9pRzf/z
fvcPWUTRaUVGMGw3OOdlCBM76itSEJiAS6lYgoL81odLNmPPvXUhJpK4OOs2mf4w
QHqFUJD2Jfz2ukzmpGhFpZM4IXQpMK1Cmyg78j6bUjuX46+75ggHcpBjShr68JZr
c2417iHiUlKylZlSksUshlnsqOXxkNM1VY2Stjg92Dq4l8z5VCNxrq/293JS7X8q
g86JrYWyVYX411jhwuw/pWytCTwtNNTaVB+YeD0SQJNSshMOhlLq0AoT38K2e1Op
0fZlD+jZbF6DVGvNax17ieFylo9B38Bs2LA6Na2ovNCEfrQQayEahFkUElPKGgHR
j+4NSsX1ztrzzh9m2s/J0hdL2bvnkCu/Q+lg+68SM+jIHRE17gw7UFE0rhbhDRkg
9GuUs0B9l3RVXu3Mf0kOXXwBNjNeN0tDpuPPbFys3iBQo0oEJ5IW0nxpQK8LSwRX
m/m9l46BzUAMRwofD5Ra/q8Nav0uhi4WBKotzwOewThJqIjlHvO57REeMORzQgIB
LY8+bso7gwXdDniPY8pFfTh45EpEebQlO6Xxnbp+y90h5G7uv+qgtoUfK1GVAiX5
WQDuWYuYURCgyDECB/oRI7wblJmZeJlucBYxzOTHdJbUVyi6bYMNisb0a2phCxUk
LMIcrYtuFO5eAWXC5KQahKIqTRUk+PRSUsD5LherPJqxXiAYvds9BUkG9/OSJTI7
ZatbH78lJ2hCdZ4Evb0KNfcHKLl+tEgEiVX0vZ0TTuwvlmXN4exHyVOzgoauWpaR
MlbcL0QCuiZuHaCGe4lXEImwgfXml9qmSaORmLN+PMaizSa74kzDILxvrPbB7RYS
L0VMt+X28dCu+ci9N4sAsVVidaj7pwrIt+E19yOT5Ip3+8ZijhDw80HJ3bD00cN2
El6Ivxccb8bi0dTFCE4j5cqaMx560Aj0Uz8nY3hIRSKUvd4hw3KAFIgNoPzLvCSS
6VkjBu2m3E7GWhSLPn9Xd7GLYEu9uiEi0pzCALqpVWcNAaAiBLl4wW6cFa9B2fOa
1ClIYXYnwPDLiIEDn0tV2YgUEUDzf1LV5S2rUA+MKFcweuI4LFrFQOs/H2XwhlDc
cezPuRMZGCORjs8oXVK/Sw4x3SlfhgvsxFasGko/UJ3QYwiHvYcL6jmHtHkZwW37
qHXCmBrIo3f1T2CJ7SAC9hW6FhRgTfTV/jZIXz189colcwcABbv1pbXRBnNin1g1
k2DxFNqDJRT9a99sHO+0HCPngyZxlXn1y0lYPkFHpH2m93RHrTgo6wp0kagGG6DF
6e5d9N37fuODTGjD/DUkUEIo8kRrFHSGLWmOCKSiY7UDmtQbcKxx5tkQdhoFQDrb
sa7IjRYQEbiUFjttxjo11e1h6tsRoKp8RuOi+QXPpXGjxSAGyag4QvU9p6YwCsWF
tn6yC0HBQ+JwXld7k5ayXMFnsNFZwrqZlojPKvmN7vR+jtu5gs46SG8P/Cea6NRB
/haFFmB3q13OBo2Jumb5N1/gxX3dOrahGznKr/Qmlsf302368krAXz/CDVM2sw+L
0Q4imhCt4MgTBWbTQdTSahzvdydrIhSUEMdwAB2iawvVn0PZvoezCZSzcP5DGplm
D37wnVXutrnmDZtFOW+HrgwScgUWviS/Ad2bk1npkig+gLx/DHtiL4nF/ngTh3Rt
7HRkBFgWJsxC3vchjAPhf6MQ9eQqnDCTeUh5J+19t1A4GSv7Of71+7M9J2vZ8beJ
cMDWPAyWdq21X5fONBGN0NVK7WTKR/HScxc6I63Yb26oqeOsHN1UcmZpdeORh/pZ
gZWLupUo4uESJdnwEYvWVi+K5zaotzuMEn6Sa51qEdtcDAQBITyL7iDxBKmsa7n3
mNBU5dViWXjmz9ks9dEGdHyjiJob0wfJbMqa0hUy2Fwv6upGl2Xi9tQrb+NyZ3/0
mn6D+zj+W6+l/6lkkmmbK7xPFLU6T/ZH2vRwOznnGdleQz6NMb4y/YKKteEvOFdl
Zso/gJ7YuJdx/F9O+qkxJFaCmRx0Gnr8SrDg137U3nETwTppZ2toSX1P9y05V5FF
iPeH4uX0/WWJ4cB52iWl4+kJRysGlXYoDui+e3EblwFlBPozDyB1yE3zHLlJjDuQ
LLwNQl/k0Mh77gGJpKw7qZfrf+q5szPEi/fBux/9q6QIDuDyL7MnKR0Iw0eA5Lk/
zZAoNZ1g1itkwDeaMT33iXelm9aWq+jUZoPjdgjrTPpMlzVzTpdhITYhqgiDJ/JI
YBGdt7aNyo1WxpL+1GKV1jNSMUKAQEUaqB8CEHS8JYnSScltigDAcLmj4ZXaFbHr
7CwVj7Wlj8S+kcESjV3t+nZCXXxlyxaUENU+XLtHYS2GEBiuerXup9DJEwjRfgHn
uU2jCUyssnGOKMaxrEzXgh7gQ6b4ma0Lb0+UpVltic8InWTL6q8X5X8eDctp2l77
bAsmrJD5Av6I9nMVa5OP8fpxWjNuqZ/33ktJbbGV4KIuSYySX4heO0rBo1lTJaBJ
uMrpFkPnfbLC5gHT5jYO2QsPJaslG/VXF5qtHVhzmxkGZ9vLbEjnlrPqAfmo3bds
t8jQj5oVRO81jb7DlTFvb/C5TWOxVxteN6PrYYhBXULfmkTSlZppHsfQXmdyZbNm
3bqrBJArZ4dX8IC04T7Yd+nhI3OERZlw26P54O1qZvlXIkvgFGwx3k7XwwGxjT90
Btmxf5GgOVGERF/mDBASzEWhd2psd4Fz3BbW3jhiQIBNErouSqUqBhtCA/D0DQFb
68tke/dATtaP2a75dIm9T9YyGGWDZI2uhmMp0hIphcSp766hwRW9F597QHWwN2A4
SOIhaZjCNhM/g16utfgureZ8LLkr11CwVJdjtZNJeFfjADWzHkh/mc/qYnB7zrfT
D88TMXCLa54lv8sRFtM9Q2LHWcKr2Trdc+KRcRpSher9F1IENSNYUh8S7p1CSlaK
v7Frr013y+d0qBDCtN/+EjLHPDzS4MP64w1+kp4dNSM2Nhr/06C1wnQVUtkvWyQS
DCg3GdKQkMk2Ba38RlTVMqa8/UrSMImqf+uBI9CHEG+Y8pivx9ieZQblL23Gik08
W1ZJR92l5mntnNawFI+s3EynWeN4m1uY3rhBG/vk4i6106MXdgcCg6jHfhVxyCpe
cYJHWTzAr98/1WWOX7uADarJiiUyEpdq5gyoZWU8Lu1Us4ibG94+kJ6NqUVHZM4p
iBQFuOXo+yLVb5mYVRYJGJ5O94B2VZ2/TcekxbCw4x3q0V3ueIYCbTOI4528JIwE
B7Jz7lmo02PPTahFQq2PiFhApKRRtQ1LDznIPolTkSe/NO8QbrvyzTLfkYMuMzEn
vj59gbT7HzwNl4JSzr1TxQSClE9vUAvA8NH7qY7jHxWrwV9f4ZvDvzs7u+/XOEK3
f+N2P9DGNd5gopM6d10pLtvAE+AMusaFd7XzVEszN5avYBTnbmr0eKSzy2AfRwDS
yHkLSCyY1n7qZ0O+JjRGyTXKOwkH3k+I4PMS/fs+TCRj18cLHbnLTGYt4pZRZxhW
ywuQzN+OtSaNZ+dMwXYStz10yLYUQWIwmHY1E/2Y4N+tznKrklPvGXp9IwQJtILX
2KsGSgJYFK62H7tLtorNgKrS2VJXUfgYBWxJVSQWmlU8zTWF/mQtedf9KHOw3GTB
zZbERWzHVTc0M8IMl7UBnEerzq6KVja4NtyrV0ku0MKoxgHFFaHQUy6QqLv3BpZ8
XEwgCjWg+KMUjidklZuXrq3MfrY6zvzoAPXoFaY9eTsTGVseViEcsxXHzFAE3tA4
oxGuDtDN7kneFJRPgED/S8yYHrJjQUkKd2aWv2pvt/PBrfaGXeKiR2Wk8xFLUA0b
nSpj6aVOCm19AktHWf6/OYsXNNHGNMjRzO+NiQWxvt7E8OMS4lmX8LErcEsW2110
D+TXv76c16JRX7nykcmVuYvanWEVA219x/LwevDO+nNB7NLvvh/eu+xFqyiAwDsU
B+uCZX0xSuuwtxrt+MUnRx28dB8dt+qhb+GZugOsO3jmOluLPU2FrMGeNvXs+x+Z
d6hyCacYQ50NrvzMyYgFevBanW8pppF9oCTELhvrViAfhAkoTO6gsYX6pHKgecen
1KGKrv3AtusoOpUyDxzR97RrmZ+FrOmZ/MaZ7+WbCuArniiMHxL14SwjHgrpr3+5
R46hLFJbSf2O72pCaRkcMP4o7kBJoQqJEa1Ut8+dXszowVF2S8rf0IGc9h2hYoqL
SoSPa31TtkjUYAsR8kp+TOZ9Dou8fwfblIBuiea2/YdF5Nw/7HhbfzRjghw+ddbs
XKle5/6qDvQA9KyLe+1Q9/vdv/VgGK89AO5UMmRiOBLWEaWMUb81IeXW6c2+2VHR
cIZQR6lZy2I007jDuxyNLTzalw8bTVPXKIFPbmkeCxD4xGCv6UPeXOXWlSuXMtoK
8hquHB9nWsTnOGOXTZDgvINQtOVKs1rEmbp6DgCulxR12DkAuAdSqmxPmJHhCgAp
kQB+5qE5wy+RRvjrzlZwxAz+ROXP/DrMx7lG1KxIY94XiUqchSmiDlfxd6Sm/3+m
0atKrCHEJgMcL6pgLTfqCmmRx3LQXcfj2WnJ6e/doS+MsR4tbBZ92PhU8DynAqjS
qYQxhDI45oOyL/qLygOTZV22wV+trBzXhYbQCGTASID+i8MmiJphiSGL2hSbfuvi
5BxoCtnwj9eX0LFCQnMMCLa9RjI+fX911B9n4LuM5YJlHn2VGq87u9HDZhl8PNHm
mtvFUiKlDYkwHq7rgHTZ9IfUJ9076KGQ9P4TAE6LH+sNu4xX2J6vxOr4X/YENimH
pb2scPOAjp3pJ8YbGnNKNIR/xohBZ78JQqvOwoDvfiR8mtXTqbGBwD99eQw7ggue
B0A1Aif+vwFvxi6ME0tNniUXyFMRC8MuXqbmEDUxRk0vbjUhJagwkS8mXXdBBoel
jglzofygvQE/FpHneD8a6PkUZMCWbUGScLYLd68/u13qXYgvSuQMCpPThk3BVP/g
Zf3g3sIp7azuulIu22K3dHiINUCj3e2bQYf4SGKs0VeRFuSIIhZBZuuUv/2vddhZ
A7w9jJnSN7XUOhJ0Kl2aXcukpLZSqyiYdKp+A/IxgihWocgf5HdF7AWhTlPYdLmq
8EQ3Dwee5WovdAmT+DrUXCFHzBUz2i/jinlOhkebnrY5M6uKc/RK9eYhyhWiWic2
5EgR5VRWOhUtDW661rubJXe/+DkhmB1oyGe2PY3MFXj3+goayJLj3qatYQcURxwL
C32NNCa7b5BPa2vFGmocpRrK/XZimaiG3AkgT0r4mj2n/VkLw5+NsWgsJAZE4sNu
HEQktFTTWXy+4d4PynScaNeHNckUZO57Cwoge2T4UmWReQml7YOTh9becIRHQ1NO
CSsr9bq+yrldusOKxn6NYPlpP5bp1eNtYiWXiT7r0Qx5PbV6n+BP3OJpvn+64Q2Y
G4VhUoTUHdqr2RKeMvwlQ+X81G1oYIrZ9COHVj/2VYnbi9ne5Fd88YMyXGEi0s4r
mh4Xc14jAxRW2SiLqShk28DW1k1FCut6hthi7oICILdLYQYf+K4HLoODdU3JPYjU
cLr4K9g0NGN9BXIutIy4vgAmUIXJONpfWACb0NTh/BzesAPwMgSZCZUqckujVNOl
cbIPrIo9wrZZ5p1kw99wbXX+0SErRRTpw+DCGRX9cvlXXiOHqLuyOwn6uu7scnMq
Wrizo8noA3jelWdvC6rjUGmi+Ptv+QF4mOyWzLfGDnuAG6PeacXNbuOCLQCJlWvm
WloaZfYk4Flojoh9/QIPl6F05schEQUYYO+x0/C/uPaQ/3d3U7nHdZvin/BlJsFD
wNPydl2BRSLflb0OUlwAd49l4SYkMUpx5WK8ijiylC6q+m6Xn5gLYKIz4B9wQXir
SNWSjOIgyrTqdflA3l/V9Xpe6QAs1Ci4r4nShk2IDTT9WsOajl2rAvNo9wxAMQb8
YfBHR+HoEae7Z4UWpMBBaoCvOQrdcJieQ7T0sTl1yjlSjAXuBH6onmvVIrsNMwDD
0B9bnhYpZRp3llpwcz3EKacXZ1tMbFKJMvlPU7OGqLVNBNN0YuWi22BGQrj+mDZG
dhYfOB+TMHMh52grGcWcUl/Z7qE7eaIWPDhxXLyHb/Sf6RByUj5UUFGaTJ3AV5zk
pEWA43MwuICYiLAkEy7X5W1wrjyJ7CMK70pYxi8vyDvCYoNGc0amjhqcthsQG3hJ
tFXbTw1LC6k2ZF8jVgDR0EcIa5L9G1mYazzHEAU8EHEBl4DcbfXcEnP0Frq0vz/2
svrav3qXkZoa/9Z9qHiviW74PSaW1ACZny3eiIJQR7YxRhTsl6fl5aEOlizFuMGz
5iAg+JGvehKFUyTDhTg+Y4bp/Duw/MKZ/jCOFG62fM84msLziQ9jOEPsOrO4K96/
h/SbQU3rILYrZvQyzkk9e4Dshps+U9Uz8xN82X4hEBBlbhyeNy/2/qjcmEGMVzDj
xDtEOh1ljNbZCoIAwoy1Gf0RvxCvzkQCXbF0VapnSn7B7AOx1FCXTtnpmsoh3MaO
EK5hSLoZAM35L2jkD1a0jZPadHz0JIk62r96/C4tmQVvrEYaitVVRJ/CrVrlKdT8
fZC+wzj7+gXP15ku54gLfBcVoLeGbbNeiaWpXG4M7qhEsmQhQOPxBWaN/NRHgtZd
5rzcoGk2N4xzjinQXxgef41i2c/4F0BiWJQMrrAJTByVla26EA5RnFKN7LkXqDNs
gOCv/NxbY47N46Qv0pyjoUPQkncHqRQETDHdJwi68o8cXsKaFsrjyd0zqCjyhr+T
Mc6uvrAr2IDJD3UFk4ZJQ3rjH4rGhe1D86BpC9l1FUyWNEcnlq3tggpMuH+PtBjR
R7nIqzS5KavyxaiqMuX2sMGvw1OpgRn651IqRtIaB0k2EbG3OxAtNfTmnlEHCgM7
GJcRkyEVYTPIyYUs2hMdHtEoeNgyjtf7oYahkaN0XCgfJJRFDT2yIMFNlJ8i7dGx
7mvPTpwbey682zhm1Q4M3rvFaSfzPy7r5n6ztHkazGsPoE22lr9b2RPwPYSb7pkF
DtUGOi3abjnLye/NdGqoQCbjq1bozXqUxmcx/Hp0xvOG2BChjCE290ff0dCOZLIg
ItV9keQ8mh+O0cHOmowMDM6aIVqokC0XBska4voQWsZVkIEH9rAieW4rZDqmDH7z
jUmxt8Pv81kmGNUrrylBYOuDabv6vqhINOIxUxadlYnM/22YGW1Zak8BhOBjxDBX
BU8eKcC90eWFOMq47y5iKatzAEaPR5hdY8QyctJK4KZjgTJOA2Mswfv18uXP+WUi
9skhQnh6S0NaxazHPBjhxtpV25nSPOISHgzW8IuGu+hy89QNNUjTELiR5ZY/ZQtf
pjv9BXcuNRg1k2GsInNoeu84xkz4fc/V64RAXAF+7SU0bUtm2G6aH6lNJuYpe5Hh
zh4jTUn2S8A1RoCsN9WxiSDNEzBN82hvH4Z6HWrrAp5RT6DOpE1xYkTgPflzNUgy
e+CF5Atf4NJFN+lT7GIWONO1XBGQeFgA0YYCLbrX4W+c9UYRVPIjGGBoOyWTo2kg
F2yOxmclheN6eNgokVA5NLWdI9DU9Cq0ufj1o6hVPJjoDAJv0RRyqCNx60P4VKQ5
+8F/UmINL6sFCJRb04PsW/Z/9ywTIlZf/4+DoKreghTHRLdapun/m9obg5e0+aq/
fsqaoCCn6cIkEXMly/RznjAZq9Q5EwnxfitciY8FzW9YeFPvXjzFjUJXKHw6miFk
P4c/lSQCwnxD6zHdrEu+nSjWxcilMDoOhkVdEyP3p4/Co4cuRzJ8dmtqtJ0fNtZf
qsBbBiaZSoYEXMHocy9JP7+k6WVWZeVwMZ0t8c8X+a5MBKkwW1pJwTq2iUYd/rmX
j5R2cF4QhT2MuRo0Ib5WIURZr9BecY0JxMqKw3gJ9/OWRtkz5oHpGopd05OdCAqN
zEoQqbENwoDrFcVaDjTbaqVS14zvOVfAYhkjx9kIF/5d0BBnzya+KzwRc6KDJxwk
zDslGdDO3FX2IvJ3dfcIaOJ2dSsznjISBGUiG2mBVTAfkIGsqtRQhBBYdqkWMpAb
ovLENgwzTdX5OHD4PGSm3GAeftH8puorWtlVoNVUw7EGCdqlJTjwCYsZTdpBAxGU
rhRlaVVeaBB+siJlbUHuR2Tduq0nBi+hksKE/McMDcDo+ikvrXTldY3uuxpjbmsN
g0qYmr8hn3GtKv6V6sQBNWL5qJ+Uv+2DRWtDAOtUiyBiPLsGq0YKTbgC3FrtbHWa
74afNqY8/MXbnwzcLWFHvHEPi3MZJFFlqX9U2BwgOuY1wtqIhMFJ7g3lMrP3fcP9
zW/3GT0cuMpmlz/yIrj01Lr4dctf227Rryh0sfOhHh28PfQeP9zYS20jbbIljXqO
84AlbEazlnXGh8swZN+E2lD2nEMSz1wwf2TxqZXs2P+2d0PLS9Sr8oDK589fPRm/
rZDtLvwiv/J5b8AFtbHh9MrlO0eqzCOJ+/iUqNbFkrp3OTNep8UsrYZasdjMWe1p
TC3nyRnyFdQSCqGfGGgCqsUKL5Vb2bIo5pyvhrLQjWdTpSfeUDzviGklzx/Q23uY
CbSFjJE7nGmJqWLk+CGHtNbw4PU8IMQbBfjezZqExNQtDZS5c1l+ds9OjPTh1PZp
JQS2nS73p4+BGBGQst5/V6/REet02XSBCSzmcByUipcrDUwXRVzTOY0Br4/0c3sy
keWqCdedxl5ZFVaonNLlJyM9fePLTrNz9bpqzOhZw6oHpDhOGhLi1+LhQfI5yzVl
GYSx7Xg+rdAVxdz58iL3Md27FJQd5w7F0D8A+9qkxr7iGwZDrwwl9hbxozPL55o9
aa5Ex7gHVeU19k+h9Dv8bY9pkuR1cJ7JPrxpEs7AL1GHl352ETwg3oq4IYDo7hAU
L0aHmybLOpuanTkeVUU0/OWZYyuTGlON8kMKWP2EQGk3quuNQumMuXJiNB2EIlhC
qoF2PngAtyGWvczBMgSRtPKgCOW1plSGSz4pstQJDgqIJzYIyjZ6FNziNnntt8Db
NxBrzO5Jo2htpgcrGxC3rnCc0LsUcPFwxYVPYYb3Krv3QSLWdIF1UdqgTMXiZAFs
gFww2PnvHMSGJRIhtgJRk0hJ7epdoiaMFz2ytliuqvrVonf/6Rbky9XGjRAP4ipS
yIi1PBAc8XLpG6ObJI4pTiwp24xFnoG1RD/YGCMU022Ysgr4r5n4HfXBdwWTzTFb
dVZzNpLhT6Amiwc8U2sHn0eY1Bfo5xvlZLQMlWB9O/D2so5Txjc4pnXFLwt5ZQV2
QcXINY8BN3ShlQtmW+INs2mTs5A5X9DOU/LZ8bOt9U1rlfsnWvJrUz1wHuXM8rjW
RG11YfdwgoTwrUFTpvtW1mCXY0zR85R9ke9O1ADSqy5V6SXGjXX2NWOvZCizoDHe
OD4TFI/UtftDzTYU0fp3xrrUKKEE94OthtD3dw+UaVIz08+9Nt9yNjkq7oIkOedI
FpfoC9jOquaXPxRvNaxSsiP9AFxR54jH63SuUEPwF8mkXL3tZrrg2ZiuVZgbVJqT
ITfUw/9QGFiAE/G6emchXW2Lkq+h4KrTjUT9CwrEA31SGusnJ27F720MFJ7YeLMR
cAshWJxmcLptbYE/VXoE6OaVCdbFUsUDthlTwX1bDibuezLY8jysNzN58043pRl+
9xIqu9M4yLNJUQXcC5jgdDLM2D622xglNPMJxdOoqkVVHDh1bDG3pKLs9L/MJYzJ
r6MxL5SktxOpT9r8501IDCbISSMEAq/0lIlrGpI4ERjQgoeqexfdPV9Fhd2PAfxM
aGF125GSoManqjQfaIRGwWpD6LteZE5Kv/ONNduGO+BKD+s92V6s9plmvL0d4JKP
ykQ8paYW3vEu97eRxp+z3gTbfKLUuqiAQV3A1TEy64uJ8s92XzAeRL43vb7VtrGh
4fiYNq5iOJjC5sPbhVZPbT2yP7yg2Tfz+GkteIWVnm/X34RVCmjjUNA4kaOjcbGf
mtm/bCqM3PPWfPZBYjtK/OiTiX7wAZ4Za3rJdJBGz1TSQd0WOaZKhAquZ7xDk4J/
Ngn7KO9M8dEc3kBwqK7RQ6rgq/eqF2u8XAK8yLbMsX+SmZ6v5r+Gsk6KviMtz8k4
VSVSAt4vFrrzgsB/7COJlZDDLzn1hJS2syRylnhxuC3Ygu7dEmAEnbd2BXPXoore
JEilCiE2lGjZVOz6yZj2YdszU1phBgP/zf1snps91hAplktXtuZncrVETmw9jikj
P64HzpGImckdt9B9EIat0nwdksH/ZlPcTBdtoK6cJ0y41LBXN9VNzLihkVGuDvol
krHV9mYKBAYLnPnYKiE2C1A39T6v9cQMdcxmZkBZD3aobAGuHZN2tNMurbnkd7Ps
Nr36LoF97HjGOINRWGTz6pHmakwAufMy2wX7jLw5jQJyg1iy+z43tvhAKqYl+P9s
kulj8EaIPvsBAyu0xm7Md/gMNEwQiSr7Mi14z5HTOvN17jbHNSEbQOAAs1q+XYeU
5wgPXoaylCOCl053Vz+yrbT3MoiVy3344Z4MDB4QZGJ7fRXahfWBuOHj63qVH6ZG
F+rpQZDKUo9Bzj3ZjAdzFAVqwgXOCeVcKVV/bxptnKIP/xQHEHALJKyFpEKoaeay
/xCKg6Fe5Z/safxP73VpUpmZcAMKwVCJYinqB5avrqt8kqr/TaExt29xzgO+in0t
T96xb53hTzYjC8baJnHY+wm95LzPBgj12JQ7HmjtgLBPXECdSSDpG8PaK0S5Eq4K
yRUYun23mxBOjvxQmLrWp2FrmPZAbD7bIFHh3XoqOVxPFj6vzYee3Kgmn5SSSFTK
QmZMsZ3fhDR/kmzp9fggsSZ1sF68Gu5xSoDrG0m90XcftUb7jaf4GWRfo56EgKV9
DCq8rZWVsI2nboz1AkwVTuuJWZmcNocLIvHwE0ymLJzB0+4R+jChGidrlefQnyla
GkEE6hECOB3eRuMzmr4dSI3fifu3Ysk1OKGMlbk2gj/4wktOirMILxPROzZZDVg2
C4lWg02EFTebGTXjux+OgwvBPtUIbO0QggZL4xI3SyUlZCrQ6OLkGC9DKXU9GFOP
HTAtDLmKyqF/sLs4jt9nZYDrnpZBieZrC4d0+WigNdasnMY76Yj37LfPK+IhaBC+
1YdmavnqlznymFzPI5/sKWEQC51PfO4wzD63hrAptVJQ0m2yTmDJT853gSmfnhYY
p8oeTkG+9dJMDyxcz6q1gIVBBDZCR9W6lMkHh8H3wnJ13e5hWoJkgwyYvTSAR5/D
HsGSol2yQhKS3F6F7NjGjBIrQ6W9hSPrfXAzvrXB2LzYgWIUZefvKiB6qbhK6HcJ
VFpkpVv5AyvplOfZOFCNEaFGqC/gGHaqJDt1b2oKpbmxJCbt/mAsU5DNivX3Udih
fUPOdgkOWsyOSydngVpQISrgOrmBJLvs68Ylbdf59/+auV2wlMXdEprU55w4YmEC
HNjdgV1D2yVpgQNkPTrhgWWMU0f60dLiPmNFxds9m/5cJLBi4cMpjrzmU8iAn/a8
KFbceWwmyXUM7vacLBFt6P2xLl4WuRELBP6HEAOCYVqux5pwFM9sLuQ19W0oj8gV
yg9G9mGCPTsmVQQ94rDwiqWap9H5JTq8IB/aJlf9Y6hcujAanJgsulWI8B/FMZmM
8vn6dgJbdFG9uzgEJAw8GlZDaHlTZV0+wFqqFkZoCAGhJVVgssGUT8zavOIA0Rre
5VSF5cwCAUPvIxeuMjokT3qBRuNgpdwA1hWRzewH2WoZsFAJLSGZ0nJrA4vyoN5n
gwOPb4i8QYEKMbC4Fv4wHf3B7EX4Dl4PrKU50GySfgvytyrq9fwdhdqoaXeYZzyI
JpaGMPHUYgDEQo3GaD6VCdQjbReijND1l1QKQlCLDpbvSDznmVFXttaEfdBTjOC0
LJDQ/kJnWdo5xYdxuvPunr4qXGw77OnOF2Z8yBSQBVWLy1DhVDdG1GxvSlGNlfPd
/pMpzu0qwBA6X88HYbgF90XOJkPVPHgsFby9FGKhkT4WcKVv0uEu8osUUybR4RC9
NpjlyRzVCribZ6xgaJZmzZPT/AxhsxFmwjyEmX7zmDZAOp8Xp9FzaZDdUGWNwvk5
3pNN0jaZQsTJdIXNfqxpwQ+HrGZzieBsEFs++HB8l7C8G8hWQz+rFBesYkq8d2gM
Qqx6x6j5izD1Y8U27CJwEm06yuz3bBXueiXMjs4VnEi/Z1dztaBHpVtqqOydF+0c
tMwgTubyULOY6i9uUkh8FUiL9ruAK34bcrM2GtLFXaJd5VFHMMPS//IurDTIYEmJ
g8oKGmU5/V4gExFYnmWsJTNb9NCusPw1fP/Z7fMAoaBRRB3QyKNLJrUWLgct12rn
WLaZgknZvP6Fc00sX7LIt8AbELm1WkmWm7pMEbn0Is9K95V90TiJPFdGPduuWx2b
FLmnoRwfO9SXxeqxA0ztUORs/GyIQ6e2aBkiEeLB5OUNWriQxHfah4GJErk9vXie
cKpLy5gLQZW355ol9ii69RnY1k05iDKLLkPW1vtI/2tB13aJtVsvdbj1uciSTAqp
uVTqyMmnrYpxzx3BGu7cd2wCxiera/1mn8dzEy+ahYkTiZYA/HsITbfg8H/aXnwp
PXBBQ00FpXnRd+CwMz/7yUcpw2U0NpROvqEqt4O+hpEZtwNhr81LiTTbe4E3j2s1
zHmvZ0pEZBuqH0PP6MwbRoRd+OsIrE0TwL0UjYgSTmYhkjUHJFSAZy6NQaf/PLCS
LgvUsctbXE3RgjaZ7KfAYr4lH/3H4rpAWkEsKV5ur2XNBfzrxmu+qMhPCko9iwpt
udGJyIoVG9+QQfsp46i6/DY4Q3a36nAIClFctgUfgc0xcpCZkVTxOeKKt0mx7VYT
TF4oR08ll0Q5GRUCcsITh/ZYVHt7TZP+zR5E9yvZXWNLPsS4CdUGLJyZzgmqThuA
JI3GZSHHA38m3tawFzJCy+IvNAKwyC3vuRWsLmfKzKAnRvLcbzWXIq5gcfKc5r32
Iu81sj0eSXNCUOJtSOhRKXokek5KubFQ1MjuHCRaBqYIWN4LMggQVjQIgs02i5Ns
Xs5Yq9CD1mIV02zcVD9pdskoUI8Cpj2JyfmkZiDIHwC14nRGJrFm7iJK24DVxr0U
hYpAyCQ+Tk/cLFJJMckHF/newuJTGVFN99MxG/lKh3PrejZVQTsPBbVwFYEYGgfB
VtjCgebX17VNA2cobgx4rbbFfzVso3NAZ2AoPVCts2xeJ4PJzCMouoZGpLD5dDNr
bnpCH1p+QQE8GH/9MTO0jT8uDzLS4x4xBJVStZhDACd2e3N55OUMpdJNfif/jmVK
TeUTHR3uaBEVlU0xvRWB3X56KFL/alm+ZFClg9UqNjIlGIN+k1lLK12qsxc6jhKL
45w6Swz13TKdEw8kIfrHnH91BW9dAXS/GhGY4fsN9YBiuFpSVl/vWUEdLOFYlzVP
LsCojMQDRY2okD9S2XosdfnNjx5/jNZD6M8f/H38CVBh7WyAraAiF14I54qTjFUU
w21cYgPJrkblMZ7BTwluBM0zGm40VOCmyKCt2JvopRiZaixoC4LMbRIjS/GW3WXM
lK1Gtl3pMw+B4g7jnZ8WAI4g/nz3cdXnnXq/u54aD+voNq7Hx23f142Ld31wzPUK
OLv0tCKyG1HpvHBLs9XBKukiQnp0N5eCGmHrekC82IlyIgHXukB7qZJ8Vyr2N4Ki
0emGG/zrRuQMB83nCb07AAbzpJkezvPGQpR6okFufY7xvvWWaJYjzRGEoS3s2k0J
3OfAgeQ0efY4z8iSz73PItV5hEeZ6X7hHtx2snnV3ZfM602mqLP5DOITdkTis74y
0ptV+HzFC9PptQCFCdcZ++gSqPPQz7CztykstHIO/CDkUQqdBODqPMP0/I45A9Sx
Qz65wf2qd4UDkgbxDS3k1PJcpfBcRsteK/b3ogTIhBZiCNUnzFBE4CmnR+T9zXNz
l2+ovwTeoNnLo4v3OTvG+1GcVkhheZm6Mh8+lNtjLyShsgBhR6VkX6sQndLuJyjs
YvMF5P0uUVZ66BErrYpzmAkb2bd5AvD1WvH+Feq5BCsshX7nQNpBFUNdRvPoR+gd
Pd3weWLeQ0UqmhELsBwvFfQ9DvJgzliZ7BDVpllvOZGFtzs+stZxjrUxDwifQQxv
W4qZWt6deU7tMHSfdGp6KauAhgYqiY7uf6x1hdecdCud355mdHZuzUDQ52tPbZEA
Y+l0wHqcI09+1t8v9Y3vTTFYwjcrQrPjp6q+pyE7f+ydwW6SbQVf8eUYkt08FcV5
uYX3xXy8yhACfVvIyPvfp26LPT3uBp+GLtlubV5VR93VYF7mzBhCQ1h6akPbtoMd
Aml4dtwyUz+RgivelwNMKFIihKAWmt9ACBF6nox0up1AQvo8LTLc3qqKPw4UzasY
qKTKE2+PaqkXsj2UPQsYYob/UGVDZdYGPt/cJsf/okcrLtpB0UUShXWN44KeFKV8
pGwfvkW4yhraG4m3OZ5lYUz+Ieeg3I+4aJrgkCfXPbtAYJWNZPqyquh36xNV9CNW
NfUmIviJeliOo5tSzLglE1VewQkU6PKU+x7AB2vAm1fvv41k5AMFUAYmjzDgsVwc
ID3NePoq4DIndkPSQsH64lhrbFcATownYUCw90XjFQKaYPRs1toGPt64sjWHD0Sw
UU6IghYjxpOXNRGCOa0iYmBlINf2JVauJikOIIKuEnb0AIUBkPik7UrkcQ5FOR9Z
wzYd3s22DEoYpOWq95ItT9CQXTt5kCKEsEA8HXwSM6zVtWDymy1eiIhc1XrQFKiJ
jrDs1y9O6wHNES1E/xp+hCFePYcFSW+VPdsg2eHNfO/64J0IuaG9eA2RCRpwfNBq
d/GCAsIyBVdu5zP+yLvUG206C5OZbJAuMs3JcQOAEzz5+GVhW3GwJoyJpI+g2ZcN
wn/V0NHNJwkV3rgg/cgdSAA8Q3df6kLUH2t+y//hx71LuOMz7j+BSeRJnifQqtYu
NfnXDTIBssKf6llBz/KmicNJJ8Kwsiteq4sV7s26bz9Z0dLZpUI7AQ17NnUwQKG9
wmh7i0+AesNRU/IYspP9x3y+huIWpHDM1MQ7BS3LlweuqOFm04rUOqgu5MJBEEw9
jFte8qkHqKG9Iq+0Tkl+x2qQX2UuF5l1LHmy9CcjT+C/4SG0gLkPEQ/AxkK4Zwyi
+bBGPtPuP/k+4x2rc4bhGb+6WWjAHuP/+yka8NuftLp5Wxi0ufmu+wcA+7FJOhwE
TsN8UiGb+jIGnSsNcKiC5umhvNs//YC8OU01aMCHWRfgLHBhaLFYTYUydA+UH90b
1zTQPerTxFVAOCn6o9y8dpXpgvKaVapeMZTL6aRVbWvTQJBPv20MSg4uQuqMvKll
u3bPcgRKkU6BALnhzlC0m2AxlJ25bonyWrlOfUzkrOZXcfcigtLDB+mjE4ufNAKW
B18rmQ4moM+zZ5QHoTDCCsM7OCLh9JCtJognonJdmuLXytVyhIw7OgNIJGsbSyrx
tzWGXg+m4M2LV8aLYu9LWZ8cMedpFGSfP01AACwXnmlmksd7XPkeFkFTV3RzqqHw
kB8PoYnsFKA3Mm9PNlY8h0DK/fx3ZwRRPieYCbdTXFDIU/UtXO3UaFjIpIV6Afq/
cfHOizjZL+vX+DPhj+8gB9Kb5Qmn/12bpRFIwQDbU/kmwCrYtJ9UJ6fBmfYJb8q5
qldZPiGXdA7OJn2axKCYm9bD4KTsssiXLpQhOxRMuQcsIRwNPR9d2KPhteWtbeH3
VRvYFGIsqkJt/n6YS3sCYDrI7gQrHlitJ8UQIgzmP22Z1lgnjpDkL7vkznxqYTei
941askFOUKNRQlA7RIXoAvN/HM3yrd9Nn1H0fBohSHA4fHgOWvGz9u6tSjvZJ32h
X4HDVS5sj1TFN0IhHPcqruV6oulwReEFB2Gf9W4u0SsIg6og1nZu17n6rEvYxMbj
D08B0eJyjf6irXV3DLy3mIu0whT52ZPDDp/8pTtoELE8SUZk3avMweVmTWFx+ilP
OI3F0rAqdSUodMBGETi3d7HycYNHPgsnC92W2tvUq/0X3x2XM6ZoADdjSuY1cEtT
EjicPu+osQ2PuAwLQUrKMfVTEyyS70aPadlQBjf5DXUSZk1xOdMf8U+13YB5EC1X
pGXmsTyP11JCBVdMor/ltvfNB/r2x0PAASrk37U855xEs9YiP6m1xrafsyHJHAFs
QfWT3F86Yv4K/uOrxmJjOMGFnP0RMPv10KtljKqv28QSsx24vyZsiaIfxX3g8qRD
g/IVbaw3h4XVFfuEfZ0WcH6wunbyTF6TgPmV033wfdvokMBZPKVsV4HOZEmMxwTH
+msT8J0SvO5hc8LkK3swFUrmcswIwoldK1jSiW0Q8V83CYz4lTn59FEndqTe2Fvd
5vw7bpjiHRhPadtJ9OwDXfIazMQM1oNM6FTc0dLAyKAYitLJEeIOQXBNnTA9Yret
rIYpEbaMQ/gAQGnRCkM5IK5+a+8zaiyMbarVY3+uf8KVIZulbGFuS/VSpXn1xFhJ
0W22InMVmk4nyFpNRjEgsPaw+ynuahF2ruVxskg9fJPhV1ddz88318gD8AHx7FxJ
WJtFzXYQXRUEoxVAXnUuXWi4ZPOfVEjqW8SxHVBN96yEpn7GTn39lwudyo3RhnD+
LOcD4xl3/NS1khO9dVYl7fvjbhelgqG33JOIYkms1wfoY6XaDbFhkFg8ozkch5ZN
JTi4CWqEv9xeSearA/NKrtiRDwYP+89ZX/vujPIHTH6XGSWjB7a8KUCNrf3Bip8H
kav+rIC0uKVw/QeflHNvUgxUTHMOMkPTS5hf0Pa69cwZar2/YtblSRsNdxFty18I
SILWKVp2jL1E7l9mIHU3O2VK41Ro7Q5ehvKQQHScoO8KtVR6JE4OcdnTBNMB7mZ8
/PZyxgAIW65pQ8CcIXchg2Ge6tehEkUZOP4e0lrqTRa0PWmQDYvkiOmBrzkBpiUO
xf48dUxqbZY/MWQ1YKwJHiAYWTEqOQFCFCAX9g7VCqrQwEzqkORbxqLQpxl8CtXR
M0Q26WQBpUuPztTAcLdnyUOGEtMf/SNR/ppFAD9F7Fm3ptaYSWzZYJNuISXITgUB
Tp4IjOufWOcG7Ov+WVQxKrFc0lAuGi8y7yed5s1Ec9ClLkfsbT6QEG5hoETOoABH
NHwgls+JdUq/VVeR/QnxXkCOQPEK235Iu/7QFvzjnThZ7u1dxEK7D0yysAZ06Vph
+COKALku+oDhDPjRRlVCGsdQIgYlfqARZVeaTBrekyJFWDHneapZJtFyF2pGCBl2
BN3FbZdHKknPoKV72/X18+A8V+5S4schzjJTA3Pzr8Hi/GlScaJDIL8Q3OFOYTqh
w6TLZEVGtsGf6Pb2Kn22kW1Nwcna33h0tMELQkiZFSnZJ/L8SZgoorGi4U0WvVHW
fC9bAg5W4uftWH2uC2N8ozjREhW5B/vTO4kv7qHu7fcMm4jPEfqiAcf10ruXsr2m
yECGXDmA/Vvv/FP3eBlFesd8ehKas/Uv4/GS540EW6YaEoqa5FO5rizvIzhsLLYv
CTxrVrOMqLMt/vwYaQdU60ynSvuFa7ybopyM0Tn4MHPKhcHEQFNiF5Wy6megJsrH
GZlBNsP16fT9ML3ZQD08fYbYL8uMTPLiGYaYGGoFUjvIAwJ0BmfqpkCCARjEPbMu
Z7KOlFaa6eVD3+Dp5+07uffqirz5oyrDXHcgCrfIoSaDOkvIgiPSDyAAwtV3+T2M
1hg0wo6Ttonjlz9l32w9UKoYqtoS74Zq4Wg7P/IqKheGVRIl7EYfhNYmQKSIn1Us
Ail4ScJdGsIx7tq0fFqrq1CQqnAfykIr8UR9kj45h5bvffegwGAMfx7yun4nLcc1
wB2Xiaw4N2UvAJAWiedJ7uKPxkPlep/fJw238v3hqryYbhHu6Hm7IGu+8z062bsA
4YXpQ3WHE1BiAUblA9ga84bMNZDVilcgHiMpvCUw1t9DdP+BFgDZVgEiA0yRB/Qj
vrCElRuFQVYfpnbvNalII+6VKB0XoPausuNVrq0Viy4HI0C5G1yHGCZF9Vo+FS3h
ontvyNwvJwCCiEQqKvuOh27AHMkZeN5OeEKuQziy6MW5xf/q0TYYUTUVLvGWp1W5
0BDvAGru/mDjZ0w5+OEjLQ/keKqn9OBGtLSE91w8nKMAahKQDlCLkNNYnwkmUKQo
0LkT+wI0SFYN+aMFjIV31aWnqj1VTVo9VxCgYr2mokNwq+Dt7sreEzUD9pb2JGkI
aqae3OlnVZZQj1vpujZqZD2XfyYonvCmJX/NXYZuXVNd9djchrdlPYwKlUoJQ+eJ
dE1kfrZ8UbKnS37rQV1CLVOM3pJjvGyP00YbMnLF1Sae7R0NMhXoSnMpYEyd+OJs
R6n9dr9QpQ1wKUXUQ68x0MUoNdSU5qv0Q215yKBe9yWWgpsn4eOrqiSv9Hg/ATTj
aGrejojfjIuop5NtwljbgK1qaWoeFrxj4DxdvB2wPOhHq7weQ5rSv3jKjjvFXUPt
CZamT4AZXPhLntXqXqEA9FxmLkXlKtqQy8/R0KxjFXqMWMBJn5I0bE7/Uqr5v1md
kJUn+CkSC5sz8OOimi19Hr1Lamk0AwGBMSrmpCkGBhhRtH1nVp2VkIYns6YZoG0C
ZdAJOQ09Aip58ljujvTszXCKK6HZLRzcyvCnC1qq0Vyk7ZkClEVTrQBmQXkrDLsF
OPA7URzVPBl3iEESl3sJyEWPnemshAZgqCJCx+txwHM0p/7OBJIs+kqkDiMvjUrW
ehAeKiJm6Z/vTJ6/j9WDGc3rLuf2hJY4itnlfQu1mYAMt0qxtGLaoXzRzNsYsXUK
izp6OPc/Rm5fdTGga0Qt8EThdK4bS82KcXvVfV4DUVu0V2mpKnJ+4qo4c7buRdil
Q2kbV1zHbyWvfSa2wfxLJ5nkhUSyl/XZvY8Ir7ZsvZxxbHN8i3dSkkAIREipCY3m
aJNFOjfCZ1ggFK9ydEpSJTQg8ci52lU0oMtrCsNJPdE1RP8qVBZjAUSndiDlxuOA
bp6tyrTzbFdEKHMQpWV7q1NUb4ijk77qFn5pw3xHzxHP8P5iQA3BbL7GdG5U8LYu
2uoTpgZV1k7a0nPfL147xFbUyjeMXRTE7QgOkQ0Kz+IrK43QiThTKRzgcQ4ZZuG5
U1q0Me0rqvKbTMy+7kjEa8vXJh0s1UJDB/dnDO+8J9YUJVRHeSnrnlnC69s9ZsF5
6/qPeOZZS9WKZ36Ta2Ow0cVQcpQr1nQllNRsxzPcOJ4r+lIbAIjPbMSL2Bit5sQA
EGbQYCiImfU9C5SXtJ1wJkxkF9u8ko2VR7oJTw/wkSAd2jx4nP8UyLC5u8+qbN0n
kVTmCS97e/QkaMU0Vq5DwHPdkLsgNtDngvLwqpAXkW6Z2KDRIWIB6bcCVoUOOvir
d8o5+buua5CRVKnsH79YpASOjChYDN6HPuoCYJgQe1hjcCNMx2+WAl+8N9QmJRD7
KcjCka3QRIWtCFlE3/Kwd4ePZ+py6PlIsecUXFaxMAARYSdEZ6CkpEFzjoWGeAEp
pgHU/a2z0WoZgeGe+Unajyj5kTxxzGTCtJKVx6+N+ktUWANW7ktBoVfMz6bdtEX3
encTsfq3Ci6njoq8psfiH12kXH1eE5SbJpNsTeC5PMunDNoLtDKAKApsB7JDubce
XHKQnt//hviP0dTmqAYtXU3sUuNOA6HhK+VFifaZHX5jWHCb3KW0Mt0uTD+gNii2
Z1w+1h2iZnNVSVokPao89EXvYGhFDZqpZQYBIikzUUCbLo5sgPgh0NpyKS9qsDfd
YT+O0m5etuz+WRm2w/Yx1OYkOyiss+GdgjZe/l1bI1GcwoqHglooAift/uwcTTBI
KpsNiwEB0A/olz1SFKbRjgnTetapMZew1/EJ1G8VDMsIxcK6W1zIf4GWC252Gmxh
40mt+6b+7HIdviWfOre/iClTz3E8Ig82SrABqi7ELdSVoMY6u0LebHOTM25KPvYp
vti+Net37qaZ1rj0dpUUk3QeaeGGCx13dYA2sItVblAuZ/3ctlvg10BupUfraP/I
fFKNC5r35NvN6FtFMblaj78NUw/gP7LoUWB96+tvEDOjX5UvCt3FQ0d74Zph4z3f
jcARhqBbJNjLo5yZeWPEd23LUydW6DkYJDg0qtGWThdTDfPirv3nF7JzpVzLBTUf
FRFP1AGFGVq6Hm5vnUWF0v8Sco//eg4KYp1IwdzlY5QoaoPUABz6LIaM29mNRzkE
2lOT59P72GlHUBjew9n5/ccARI/6kHO7YvCLscdOse65zH7tKgf4cj+IOtHmzJQx
ertB3jNI6+QjworrlGqDN678alml/cCrSiNbY8Z8kS8FgeJfUTAfNaf9UcZiKfxv
rrHFccXPZAVI76vJmW59A7bVVVMfKFIOHz7GFRJ5ytFxdgkdGQhWDNCzpmgRhCFi
GHq/f1PfA5yM9j8v/Dr9jHNNZd+ZgzVm2VSbgIxjdh9HMxxRi6LdMTMILIaNq3Z4
hSrR1owOqh1bOcrGboT8fFkyMuj8zGMHl59IVO202iDiHj/5sxhNQlj+c7LLszYJ
bHKXjajB3pFKC5iCKaAG7OW8CTAtm2pn8IGEjCPkXfngkq4Pp9lsk+YI4sm2DsoG
jjPHoT5BARF6hH5L0IX5XuXeGPOrHTr1ITSxWuJchj07/QC4sIP+4suwu34Wf+YH
Ky0V22w5eJkYPEKPMz80k11Dq0+tHGURg66Q6alyExx6cFrA+DfkQfC1d38F1Gk/
sQ/uTvA/XLipRD1Uo8hv4DiAjyKtF42F8IhggvP+0KO0qVVeaIyPBMwiIc6OqnvH
UsS+8xo1Tga7NyFL0IY3Jj3IVdjE5lUlYRjBxOAwlm7msFVlTqljKDMt4eBPyoK/
G9gkQEoqZ1aLUUfUJ5VVHIKB9acFxWUIRQJcWzEAStU3HnqufSa5DaCwtFdNz92M
WhnEqnMo+KBrIjyAP8Rbe1N++13f3Lf6SzG3O9630LCwkglbBzlEjjuVR6YXOW8V
QUWUbOuKbfWwli8yOk6y+DVyvJgA9d5scMiuC4m1zr68LlF1hdElQpSy3ZDxzq/I
gspRQsGq68Q5+wX4eq8d0NY/hO9pqHL4OOFQdT3HYQ5OPV0h/YCSVytln40Nil1+
hGdbiQLeTdmQ3pJ8PPhYBSUgkZODcF7hH3zjI7e/5IWip9d4Mok3DXVYL1/1si+3
0xsSIkDNrxItuZqPvZiO7Gd2LqBvkzvcXoT8g6t5wcKATg5D74vVAF3vIjSVjBGz
6Gojmf7I2br9eKsNxHusIXb/CrX+nicDX0HWQZY7CN0Vm19qDUPl0SiraM3oIjyO
/0FmCnMv+2v91SgqQHMGxxf7L0D0tzUbK7Fb930Z7mWN4quhoZKA7uJgvcDDAN3m
xtCIJmQd2RC24yw7FftcCqqigZDIvr+iK1KX72oKfqAoZy0lQ7+X0a249CpKSdsJ
Ae0HM2gtyuW7cmoGxt3Iu5kYmXceWZ8HgBTLkUazaJa+O8Mwl3Qa3+/InZfZprEa
z7bkfP/Y9WKGz4Hl+f6as0/RECa5aEAwJn4O8+qmwoVGOK8gWr0WOQ4XT1hKLb9b
cyj5iH3qPBBLSfqTQ7bdJn6nHhosxolWwNUd7FjUcIZbii6fZDfQyacQMgjRu5Hc
dK1zT7zDtUDjYk5TRPbbogd8OUVoXgy+6gHg40+BzclR/LB6YGEzugAG64a3Z7EN
mv7uqhzFcfIJoAFN+eDAu12JnknqXXoawyHA+/rXfQuiKG3hvtZQAKV9taEtudZk
DfyzOqdTh+xeTqirVIgtGaBIGQDnjQneNl8tk0S7HMFbhrq6/z0u3gK4WyVQ7MGO
1JgisNfR2VzOTEsnVX048WoLPwHZjPCj8Vakdjhn8gXQPOic9+ZllxKgp6OOW4Y7
qpqMISAzh4NVDGZDEAjK2FBC3YqPSHhAIeLCBlzoDZTwq+2Vas+XaQKgEngF8Kmc
u4+3+9F29KjvZ0ZuaQOQ1pMAgHYz2gprnfPLF96t3A+xR4KBElcfKxBOybByOtVl
aEVFF+b/ofUbaZDYMA5nCADC7/D2WvFrEPfjrAHwYYhACAikoOZ3Dga8DTheRspH
vDHdGdF2fJTD/beGjBZrxA8HyeLehfX0w7u1Q84WQajXSkfKHbzKPKyUBzAlzZCr
yX1+Y0ZFt/x/+lxyCWLNCtmv59OLm+NXloxHrMKW+Mp9Fe/nADKDbIY56rembgWp
hJdvALaCxpU1yPyJH8/Z5PnhTswP9SJyKeKdjrCmaShdXiNO2cghfLEaO/60GrSx
GLXSv/1b+qaUXXJeVsm+TPjSK594fAuey1zSyM25TPOliqZ1wcEr6+1jWWkr4l3M
R+iSUSgf1A8xHIPfhJ6ylDRmqd1j24e570inNWPaZEurG1b3J8QV6Y3Gb30qOdup
qom1tov6oZvZ+iEduDb32nr8DmpvRgcRkAWqX8Yy6pf5bKOd91pqBLy1CldTjIFw
g8dfl8UYilHwUL4+e/muL1nZtxqu656Tj5ArnhtpyAtaSG88PS0Hs/0mGOp188A6
yjGUSulV/hov6xzrIw+YuXBV0kJEKTIipdCmfLM13L4dEE+wopBXFuQhC+0UR6+j
SPRZdLFb6gSM8O3svMCRlbwhXWk9XNDO8OSuB9+MYzGW7z2BIrLZX/w4THUD6wCS
zx0rQlnEriXEpEnIYzPJutzUax6ecRcwpkITIKld+nRmUzaBcsMfe7oi+XDYApI0
yAVLQaP/cj7ZuLgF4o0nznEBmy3nI3w1Gq2mPnvmzPZvnwZngeLEm+9a8inXprSx
Fhf76m2XfbemRP8edjiOVCwioY7mNB6ztHpK2B2VO7OnU0YEXGtjiQIvTQEWMdw+
nsuwhCOwFTY/0nDijmAnCK86JmsOU93IGzJH5hyxM7DZ4DVFuVzjgXaVHMor/8y3
TKOjRdHCXIKi8Cnnb6Go6jz6AcDcNwjeWZ2/HAx7GgmuFer1v8XAzjWGjvS6Kqjn
yxG1jTa1iv6K27psyqFY3Xr9giImiBgN6jHrgEHC11mIfwyBn1VcxilQ4UyX4rsS
xOxbGCMk+BZvOcVYdMKCEy/HgyC7Y4SeBFzBZxDnlpkmgYyml90SoXTrz+HSy78l
kOWBZiXC5u6dtxK+BQ807HVvrl0ocI4uBcCdSt4SKphql9LF60AG7fkwovXltFF0
7rCRwFGhxsO9JwgTDnWjCDf8tzUdm6MS6zNetwBp88MFpMxReTo4BG8X/PU+6aY8
Etj9CbrE7SCo9KtX4bfbhr6ZU8ymrIgZJdkMUD0qHludZD9lD5wjSKhXREQYiSzx
HsR9x6s7wc19Oyrr93rLZiFtt/yUZcNbxl6969vo5qaxwRD61oO/cpe9Cxt1yBEL
Vm/QyYXjKNBUt97Wlecjh38arYMr51l+PQaylK22rstu+7/uWUatEEpp+XKFTHkH
Wpz8Z/mkk9Sc32CS+qF71d7sNWveNxCLPAT8ylC7wEs9FsN0KHkmafnhuzT5QmeQ
zKWlJ1Febu/IYB1oZq/SsXynBXkUpRqJ09GOMOqmwZdMrPPjh1INyi50bYXB5zs9
e7KQm/WQtGmXaDNU1tjLZPgKWWu60BNKPd3ts+yZE+3vijiPIiirmnESKJnqLxQl
VVRejYF5uU1qGPmm7JOZP0pGKaaYHP8KEt44O0GdYajhvr+PCIf5kDMlvWQfdnH2
RZKKolyJFuwpgLGmCC2WMtlrz2IPKkoAdpkdQRYokWeIDdreSqBXDT1AhstvFcY/
Iq/hPjuw5aSrvsBLFicYJfOgzZiUv8l0szyvdF5ccR+N+aF0tDDrZzgQcD6CwSbG
kQGRMQeocSwFDnvS4nyWdWp0Qyx4AZ9oSyYZjlU3eIpPAn53irakFdiQGj9iv5dh
ZsQ4Jr7LS/+Ai63VRIa+c1SdF81+UPs19mwXn89gdAB36ATbt4NRd7uL0OCafCzm
mhOzfJrCV9OBxwds4SnmC8kBxfzC8V1Pravw8FF6TfXpt+eNm87v7fgoHSzT7art
E07GyLzm6S09KXDIM5XfI5Uan9t9rihwTadVNS/6DczlNkJ4WrDyEI4v5BR69EQZ
501wu5rjZqY8y/EKaz7dgUjPf0AKJkLBSC8CXpUbmbBucoSWCpZbTl39Xj0/Lb5U
osEwISvQfeH0uTn7K8lUrIbCW2ER3Bhtqqwmn3k6DagqTla5ZdndvUSxRu8IWrqD
8+kaIRo1ln0m3YH+GFQTTCWgahKnHDDbYZW3E/yThlFEEOC0v4b4n5+XZf3/iBt6
+BtV25i0nrMFwjve2AE85XVKBC1OazhYcp4TEuYoOEjS4lOLX4Eh6i+8bWggWIeV
ps+TZWvSEtL+Zz14O13dMJkv11oXuL1rrijRi7HFXeP5cnnJQWW4fW4r31yv4Qhz
rcEf62pfYWpEZkJ303/f+cz2hjoUy5x5nU2Z/c0ytzuTnEflZjFxwVU/l4D72wZR
Q/SMSWPHsNGtte2n373JpfdeyC0a7RVsVNh5RqDng8WC31UYlO/RPMahpK2cRoes
fYhs1NHnrPzvKub6NLYgZhUlYQSeqWJ5aSUCPOcFzxxHc1MrBvpt+mlIK6Clxy+S
QVOeXfsaA+qKFTjzvhmUFhEFU9mJ0pGznhX4TN8uwLeVC8ZPZiuJikPgmdFiedLp
kUY105Bl3JDMHbNDDg4XT9/qmszFvw9FAowjZ4CK68WAWG1lJYMq3tjwuWCN7nlw
uS9qGUr5izOOZd/pjiBqTsYsNxxXK8NZOLkXwv8rbiuuAKv2//uFkjEOkt+lCnDc
YyyqX5tm6ISHvqKsIGSFl4PVYmbE8Fk53En4ickIqDUEy+OdrSPnqAnmAx8Hn2im
2h7/1SpADSSw9Ky8swauGNftq19RjoEsSeC0tbx9U/itNafqucYNWnrDLu70UWbK
QOlWYoE59OsB2fAF09q/B7gBAby5eLKymW8zYbMbF+9F8RI+MDVyy/XxuJAjHKU+
IaiaFMZY5J+pNinNlumfPOyy/I03T4IAx+usTddrRgp47PJexLyDcwglvxB1QslH
9OQAq4S4gCgUkTTRR8UCtygcxO5eXsSqRFrNPy36YtbrP2iRFRvu8SV9HboEhwEV
g3Kzy8VmpfnE2xVCKunCxMN1w8Al44S2/CbYsZGDwkxWiFxtFhBKS0jkVl/fY4HB
3/pKd8O0JBfPyNSF2iSx7u4DNFsMHUb+TxF5UydezfLh2QA8YWL8eLb5o3TSYWxU
iN/8BYjkR4gz3XBpIfcLMJnf6Say65yPATPXJqgSeVAWZ2j8wsGqiuJowEeKuiQL
IHzF+YxnaxjqCLMDyiab9SpN3GDXGwF1joOB5f2k22bVG3dGxQf5mDwr2bEQ4Ktl
BNX3nGQFjEuWwUhHV4wnPeHs79a6lCWc237KyiLfOkj5Y9ZBK6rB8B5JFa6Fq0q7
N7kcFJVQVA63GKFTU0QoJabz026JOmRYyqDs49B+H6/KM++LnTVlRXxe1MYYnpmc
gn+kMA8QlILrw2YW3dTB95Vk1CQO47RMACIGbnLb/nFLBn7M99l/orh8DpovjY6L
34QeEvUo3sfqdrMbNYGkoyk1jC+XhCtoYKOoTgHfEp9ykF+M3+9IBXNQU61hocbm
dXydWq26iMuKkFleOtkbviG7exCRz+KTDdlvNCMU+QSGRqCagjwjclpPGusNwgKt
Iy1aLSuPbw7aJtSuE2i/JkfQJ2f0zi2ZpFZqpu4xMprx0kc7W9KWOGoRJBWWr9UB
cu7cIEDKsOVsBfZllj2+fissgEzdifvDhmZtIxqZ3O0VvI32x2KnrPfJHQHonMkR
4pz9tztvezBgCg+wLQCGx01R+/t1bCRp17VzMT4gbRAccKCwMy4KJ01JaVIdW9Vw
hs2Q+VyC8V/Mjjmazh0PeYz8HaSSnwrn7RR78V41OJdH8mCJWWWhBnHz/xJCoKwb
dK4VPzmMPm+iS5CQlxzu41CCn9GuxeHo0b/h1/1ANAaqJX9AVRXslqUR490ek1cv
9pzmm6bHinD6z/lmzdtcTv6pEimBSYL9mA+ygOv59t7VhnZXCdQ/nQo2PwstJd3s
W7l3NOVY9vOqmdNM56Nfc+oA1vdJwh5muzaBLBhyVzycHkV3q0AdAyY69XTz8QlB
1U742iaTBRfjSyoT3r2i9rlStS+w4nIFmdYbtJS9m3YX5jhzZs7E7157aSlSs3C6
irbqwzUARZumw5vvYigktUO3ZiNdnTHTVmkSNfKiMxX4MYNaP3z/mthZOEpyAzdR
1Q2qKtFSLG3l3EEks+MKaalfaWmp0wxov2fvTr6FLJBrawTeT2V0zC3Rzho0yMsh
R63tSQ3jHsU6LcpQYtgfIKAv1CAqdzJl+TS6EI5rVznrzwC0ZrZdQnD81RclaFBf
0cEOehSBKFv4NToQZl/FQhpvnxriSuDU+J7gNiZWsVtxcJuROHL2Qpq60bR/xS4Y
Xpz2AWQXuNRqsJNHthQKKMHdKTMyBrlm2qKJqXV+qkdQugehe5MefQnYixbWLexS
hhLYdDyqtbGeXnrACZ0E7OfeaHeEHFcbBfe+hc+/DfhaULjNqyvKXEk4K0caDRbi
cFsBqeM6UUL/SLYC7wjDKSunZbNp5JXF2hJ4PsZ5unGf9Xut2AqRx7otUgoVmDeD
hn2bR4BY2HA6FwYO241WiWjlFpLaM1UzAzjlbfnyBli1jCHyQ/WrTGe5uXN0e6Wn
LKKBysYcnqXaXos/t4o8UroTiwMs3tXaovBurvBClmiKlapuuWdfKmd2W9OPCC81
1axJ14CRa9JfgX/wcUH7YH62qtdTaNYy/qoGk9e4dMqvtEV1Poz7yWJNIXN4iYpW
uL3XcsVJqHCgtwmL2+/yjKx/TWD68vL4KZabMVsaHMdUz0P4Y8jU8O+9PMP0qYAb
uvHbVK7zQZGjvHUcpxS/ytrRXVvQ/hFUcx0ui8wEKvMhFuTvyreMlBS0evCX5Y2J
u775Dp+aJVrl8xvWmK9zfbE2tcji8POmiJ+QG5pA8gMLz2CjMlFJO/HSO8kwQokR
Rnx2lbC0joBDTX7TyKYov7YDr3MAtmRnMuF932H/6xKqSdQvbVbRU4wouY6delfc
DThuP1RR8J91CoRJUrhOpXnFWFCiYoYiWJA974DhVpnBh0DCJQf23c4RMqaBr7zE
ylpPhqC89tG+F+3u65piJVbGRa8HpuI/oh0zm83YSGj2SzVjl7rXNzfXJRZwhFZj
ffrZz3QtfNUdA5xJfLHEMseIqQjV6Wz41hzlfpGYGRzJPf0OTLf9U3Cm7XmIftLJ
u9kK+UAM3+WdrpPFEFUoeWFjUOxwry5uOwkYFGmHG1nR0IVg1Big8IzKA5iN9Es4
y907RZ1AfwgZ31ZK/mI6WkvQEmNp16qKmKhGrbFgRAiVN43cnPPjwPk1H2keLC4r
RC28Djuu5+NIe3DbdP/rtTOKmwX5gVrhxdQsMvkwFYOb/eiwDwrwdZaRwtBNW2o1
u92izumyTtIPLysXvLkvAfwNwOwCfVJSovM7Tl5pxuZnwLbS3nxNRLEfue0sP1+c
zCcN9p4hv5crQg6kCA19UIs54H6TSm01Esw1BgSQsB7sQ2jKo9Y0tnLN+sXvQYKP
vCnNZjmtge1HNzDiiXHINj3H55RSMElRxMwdYgOlSRsWi9gK6/KN+EEEqPxHnHEW
/bqy3b2FSy3XhFu1e50GHtElz0M+jwqZYXcCOaIt1kgKyYpIlRnwh+S1+KaJ0nAe
3adeVmP896IgOd1FxyloEHCEm+o2DEs7JiGzWBWX/PF2GuHcn0U44UjG24aNgKDN
i0OeUqKTaJBiYx9sBvDbXDUmJ3ZVtDKMijvPVOhq4DbHDOiswCiUJ9kMZZ0tXaXV
sjFbqTZXh+Qc/qw+MsABVRg1OYwr1l14wRUzzSIU+FRVsnTgO5udhcYNmUbOYrag
/9cgIrWfk0APQGgJ28156oGfGTx9IcEgdW4QXbEdOXuPD9MRfksDCP+ADRFTI7NO
FTD8ypKlwDIfe5GsECoucbuGwCiXpbAVegt2mL03mJBi6UfPKGWWpOYE943jcBE9
RZ9HDXycQ2Im3HKL5Gr5mENFyeKT/kcA7Aif1fgwQm87+EnIOYSMxqCb+Wwiwhl6
z384d5I0iJQPL7GxZBLcBa+t6cAlwdvoF9QX9gBx80peZLkFtCmtfoMBK6A41m7H
gEWbxZjnLSBc+TRqkDU3h/M6W8bBSL0aVGFvdBNz2l7tO33MUCPT7rDuD8A9ylw/
rtKl/akhsFWtBHtNOqHopXehQyJNl++6daVWDSQskHca/2h7xzO2k11QwxBCb5it
PFFddLiy34uBpSkrNU2v++gcsifj0ZIVIx6ZByVxhSbYRSe6c2K8lG3wsbszxzou
wlFXD+pr7Oy0Zpjk4DJNSR2uGCkTOvFFATXsvadXB300aXtsn4Hl6QWtK3sd84Ni
KcMz02d2MFN5wyIQlsaCmlN8hTdKSpQAX5Cqn/SkagV8/0ba7SROmgsde+AAKrJt
7lTbze2tgfIj3epIIq3/x8Tv+r8rMKPIspZHYWvcUISMQDz1FlGJhs0eAMXkdA+G
kOTfOLyGejTvIqYJ2hBr3/HPEJIDGonG7qB6b9lLxSvH/aMFGO2wrUf07PrG8+rI
ZlHTLxaePpYuEp886+fOVQupdk9ereQWl621Mdu8bB8MMJkxXXKOH2lIfgnE1dEG
tI7eHhSSF9SNahFOXxZmJUdXghhzSyYzs5Sa6n6K2MGnIatJq3YoOuh70osRu8B8
dO6v/tfkDPKsNOifb/QqV44BofKanB+mVkwcnAxZQYWrcHcjG/RHDRaThDugb/3y
f+M9IviAJ0tMn4cZqZl1sAd81Mo/TIKwmXeq/UMsKCTXVj+Q9AU1JlbHyLQm1oNO
NrdHQ2bkr89HvzeDdAuRUNlq/24iA+jUFJJeb8S0Iw55U0HeR5jqpKpELzBzhJlW
RXF1m1w53SLShKjnej0POSyq0DVnqd4PVkisuLsjNMbG8RnugyjNLvoE+ZtOfA4Y
IQX92cYwF5hnftyyGJQH6fedWQgFCQXES4UBO9njZHScG4oD+1j0B5dHvPNSeOJA
P49JRrGMrRGHl5szGfyUEZs6U2GNCqFA98zIRtXMCCUCuzU81Nc+yeG5C34JQVnd
2jQWUr8LibkLFV+bkuDI0BcTYZC8u9Pv1qDi2YBMcmAzm0D3Hm9+WI3tQEBjzREg
xbLorPtHgAMPzTeGpMPSMvPBJfVQM1y5RomLOdpWER7Vfss7huGkrc15apkQ3FIM
tT3P5oeTZikhdq+6eNuWn/PWVQIf6kay6zn/cmw+grZRk+nF+UMPD/KMBP45TsHH
89NqSJ51xAwLEn8vgvTJNsYGkla7KNZIWFCG/fhOh5X00ams7IdTYEJrD9cIy0gC
Q9ZyYHOEki0cbl81M6ICoKip0QvLCs7t6b5XJ/WhxyUJ9cyz8r4kFhrVL2XUAPkc
bEjWnpGghwpc45dx2KQmIrMueadRrTNcCyzzadf5hvplhBGSkMD1g/96fkVhnR+q
rRdsjCMdHjW7SiR5b2d7cF/HTWTBMuhKHYIpb32gGdAxQAsAw2AKiuwWlORJbfDH
DX+IxRuHKeSprxNa8D6WChqSlS/HHF4dD1yd3iU0D6KyFahqLwJt+EgEUwyX7n2O
mTNrcr3C/YMa5m2oi/OzM6eoSr++MtKsZL6VWcT3F4XVPbdhlWpSkhcIudjBoPbt
lS3APp0N0ZaDQpyeudipN2cXq66/6cV/KeBh5gGDN5Hu/AON9cdnk2RNNcNhcgG4
SmRrWNA7Z+O7VKmIBjHj+GA2nIx8HTngRlqJll02enGERBI5A++/0SBMuv6jhRvC
HkpGDCnPCsDizkixaEJ984z0gZyrD7viFFsdETapb9BwXk0EOip1ZTn8wRiRAJb1
nISpgrCdwTlONu/w7+SfJhr0WKVzv79T0gKg00VqLEIcgLxO53XSFBuXAiCf1iKu
lqhU2pGOqpPInL/EbAbll2Tn1gsYhJyDtx2TUTUSc4L4Tz2vSuj1yyjyKDlpNZfz
6ucM7Qjjj2QP4djEsdq6A4EgeqQmoqNqDPyLAjCpu+dLICnGqVGdKfTeYzbuoAuN
bq3j44NfHBOgrDNC7zknqpuWOb4HdHGTKDDCspVZ0ZxEHCOQ+/uNAMhPgKfSHbW7
JcBHnmbcDP/VkQaxxtL1pC8lPbGleOkkmMaiVGDCL+8uKUO30ddSUf9QGifF+Bkh
bhj2OJGEn5cdQ+nf3wI+SVSuGitsNKtB2cJF19Ny7jFpKpPxUHQEF5OFowO5jKLZ
oo9bEQxZziy3tnlAK60ZohldjvXR/WJ4IeJv0R7qX3h1hWq13SlrXUKpDC93fc2s
xWu7SLIl5kXoqVEG6dTX7aQF/kCmN7LrG7LqiJrvn7wW66EJ7lSkSTF04dLff2ol
dA2NKz4euMoGaNbkGRQSV25d+HTkZUW1B7hZF54qClANkHT4wSNOP01MDzAU1UR6
DAEjlskfM3efHmaOwKWLzc/XXcj1gA/kq3pu1VUTeRhUUpo3I6vESBTcUd3u9nzp
SYltrg9obzoHj4pgFVnymRP3dUO8aBcnP/7zl5k/v2QnOJOIzweYqas6OM6ilETV
enb13n51ifwSogfISsiP2kszXE7VBsEGklYSjCupAP28ddULSZKD2qCYnt99u/ki
Z48FcR2CRp76903HFozecCOKtkBaTp2zAiSjMPn6cD+60Uq0iS7COGUsISLXI1nQ
x5JvbO5snx2yRp64jOuwjSHHfdf5vV/V2k5jyMGN/aeAwP4WcR+YSHjGr7S3WOXM
y2Lw/n5rqU43mTZ+kLmxJ8Bl0sAsb/ODa69B0RmClg+PstcEW8+zQqsml+I3a+Yc
0m9+QhbdEbLbMA+9zVtMvXPohDkr9S4YfYo+Zn7L4yKX2ZYwI96VXZK/7w9fSjmN
Y0ckf3Nxf8+bfUSI0oHc7qWdGgUiNlt3kIx2kj5Ck/NMBtbwo8+ox7L9snbKVm6z
0GpvxtZXP8D1XyilIXImpCri5ArNrFCMKZ754iDCZmYrWDSF/S5PGpmaWnQzeOj8
ac34ySE+sGdwNldN/HqQa6bOo9EHeddMqlipP7epEsSlZBmUUV/XXNQrtXC6l6nv
ZpRoWS3Lg5K99XRjazB3iOXJR982L0T8KFFLKqATytJBN16ZI/OUw1mHVoe6LvY4
9vBPXXB3eEt0XWQr4aZcvQJR/VpP3hdnPWn/UTovmcSPZnplrOI57Xc9hIih+uB3
Hz7pew8JMyqgLJHMCJ7UcxyCP1yLayHB6uu0AdI4D9mSlm8gBOkDx2RAzGLn0Mxr
vZEHhXAlh5sTMdVfVzDKa6VahwTdffIrsucsqkCZrIZwu6YyxTLtfSbT+g0cn+lD
2nL1U/WRjooh9qKj+ZayxSxUaecyiNLQFgz+CEqIZt9jCWqsxWT1cwRBSSBFCYI2
O2oKuNGq5l5Bi7lKndXuSjFCjBcU9gkR7YXEYKh/aY3VbTOqc4gEDzecEAMLrVOk
XRBWe67yTAkhHfyOyF42HladGc8+uFyVQVujLUj+Gfwxu2SKUnlc3zssLVS55Qmg
bSnFnvMRqnWl9Yg18mRUoYtGIUqP8bLPzZ4I8Zo5wSL7VYAoXA2L46HDuL20hIgo
IjxBnCHJA3Rfm/HNM8KWu6xQrTP9VGPqMbiOa2kTRnwo7buOdPdVY/S0QTwIdl47
dLPEfNqr3CNZILzv+V3lOvNRNzK6jXmUHSLoVTFYWz5SsHXVzNy4zfnk7ALoeysO
N0NUqVB9iO2Z/zv5dWLES3tXntvV60yFDmXQeHiBXyb81iImOEIwC0xIYu3Aq8fD
mBpVZ4ka6VnLFRdcsyUPL3Yj22cETYJYpcBjrqcHb4xwNSZoZInWZIhcDeeVOrbL
rLkvzsl7Nv7fOehcEDETVTynDZERR1pXrB3/13YkulOXa0MHx1dCIqS2lpa47bWM
5Xm4iJgSfYLkho/FvugetzNVSci4cuOKn6SBRGv6ssm08p6T57eFCMVyHGEQD2p/
uOSZc5iZxH2dVBfH4jlWj4Gsbf44c4oc5j5fAaQi37SCFnGiNqEGczpKQYK3FeuO
bQrQ44YqNXZGT4zvrjjE4CNLpjdr6aGIr7Vj5ctVECWutGf/Kol3RysbKBt493dQ
iARbbgw7isq7tJG/c/UUgJ5qAIbp03yElfcVzsX44O9YmRLWNdMe1rgBv5lwt7u7
Pq4hcNO6N81AbTcqbGTMX2AtZHIXh5X0L9t4B1u+qYOZ+lhQG9O+rC5dTKkX4ToM
KkIyrBhiE4Bp7fI30LifdvCz1UTly7NA8PVH6o5qIeS74nTEvJZ7HLcR+eGZ8CWL
rCVpOI9ytip7lw1xXC0bVk6DA2k8ee/tzKUQL48ioAnPBuru0gaOhASTSBiQ1TLt
q+9ZRb0PaQaooMVby5Qy3y9rwvrWvUvU8u6i1cS/b5B7isHDsjs7ZP+jmmSNQf0q
JTgxPRroTpf6/tA3zimCW6UEgcIoBlV0mS3CBW128cfuujAVYlVEpcfAlK/CnQCl
WS5cWEBTvYnGxXx39Ds0DjYcj7XuMuycV21f1lnU/uGQ8ihaps+SCkvdI6wJHwFM
zfG5jqyMv18DeuBmZu+ikKw4d6IjpNjpTr/hwVw38gtenyBSmDUQGkSRuZhDP4fK
tS2ux71WNVoXJE8NiSNZEdQPJ68AuU4tOgr6Fz1TOfuYxsVXrh95K6CDdn9UptFs
TsLKaTVhyjcqzgYK6MYmJ87jxtSKWiCE92apeD1b5lTV/2bgTyuiOmV14ZXNllwC
dKibUR5NOphlQ6iTg7c3s0iuuaar+oEOw9yVs9wWwY/FvcGmzM0+UneDGqaHH/FG
ffcaX02uR521erU+qqzG4bYHc1kgSDezHVmVjcSZAk/HpUhlJquaB+vK7Ox8Gca7
K4+t4UloATB3aU/bJGAuIAkDJlP4z2yoxboon9kcTKS2phq/k+NQx+sMt5ILs8mg
T56+gJozIS0a5DPxy5/kk2/ni+SQ4DyRzBjS2fNKy2AyED0uZZsoX6F/MRJGqiy+
HMFcLYdJ06kIPGInt7gDMJ6F1WE/pGsgTr3iemPB49vcbgL3FtE1lXap2I2LRA8P
zI5Dg9YmKSaYu+ek5n/Qrlpz+tgWU1O9ZNlrhz38v2nYFwJNiPWen/gEBmZTiiX9
PsnjeNtoa7VwlZx4awBuRbPaK/97zWmBZOmyJXEPMpOQvMerpnhlqY/ln0NNjiAf
uNzjMxOK3onq55G4Yti81KCJwgQ+UiQlHL2/fu21TCG2wIzxlJ6uIZqjjBD4KuhM
R0Fs9/kXGpVOS1UxcaL8YQHI5TWBFJa23SRUENB8tlOnYW/o2NFJr5razuhEsqc6
S0GqGGMMFfMZhar44pObZ+t1V2w/Bii2mM3cv9nRh0BjMPOayWNz6MqRFKccsol+
03JeV6F9UYT5H1K71aR02bnrEm9Py0q6jPArQYkL2eKksnoopffz85A9nJhLrzCA
0D6nMcyw2zgOPY161GFQFTW2GT/ibAB0AA70YoF3hl/s18IFAxBGTilwSAD4ms1x
n49Nh6OsNfEpqa63AQriWpffo8REHwzyCwIle4IMzzshml9UPWwb9fKTYebqCWex
E7I8K1lCtKUXG+fHCvHfOPF8ui0425YoJ7zglBKfCj7YqSvBLL87RtQ8AeoMt4Qo
TE7WJO3W6vzjBrs9/tynmtLPDf39H1I9x9XbDmrf4QQqSX/qiB/w+0E9JuREvYqI
2/zKbHjc0aMROJfTskfDaxbwQjF30XnduTW51BIEptQVWOFdl5pOnxjZYawDhHm8
mllY+JTWppckXlyoNMUat5VhxhVX980/WWU3DmSvlo/rEaHltCBAEKKHCywyDACp
L010EDPp1pDwbRsnUDwk/S1Q5KUX65yEDt19uWz/uwUoRAwMiXGAo3SIrJVmmG/u
ZqAGfaomThm/O3YywkOPHk8mXoZocVK1IX7dfVFA2Frz8eZ2D+uEqo7swkxNYzqe
Yc1r/SuwHk1ARO24S0Ly9g9pcnj4bnj0XwH3Sxg5N683hlmnxPmNPxQ0SwcsvEkd
Kx/0hCMIf/aby+866fRtuIEY+McjYdQ5ZZfP47nByW124457jAHxELNYLUXRyPdJ
fWJ2gNp59Gnzw4DTjsOA7XBwkYNrICjJl819rHKnFP4mNW7EiMb6slbBXP7jePER
mOZAJdu/PhIdZNiTca5RhUI2b7s4fQD/Y80Rd0mdPos5MA+izMOzX3wDoYG/4Xaz
HcuwCfvORvEnuq6Bwc0CE3fYXItM5NZTHrkVo2vmH46Wi/hgMqagu+2T+L2Jg3lM
ueSy7meMIDYl7WBWpkeupGM1nYTIHVpEOSqIzBVjktpzAHr0Y44Jv6z3tfWrIHYL
g+NCQu93ZrAYLHtEHF/7RyQpUkc65/ox3niIQ+Y7KMe9t5znfZQM7eqvASQ4wxZh
Bw3QpOQ/5Iq03dGMR3/FrYmWh2RzIlTLeMWnlymwgtu+1wFzWo4KJ278BTTOIoHH
ejfVVCtH3AnH9x/PwoOB95XY4uUtkuNtk11ASMp6Eqv4CiR6M8TF7UYTj0cse/K/
iA0uvYk/fbnjY2J0vv137gs8ucCj5PIOXcyCPcNN2IQUdO3qmEBWinmQJWmalLCC
0ZKshReGu1G/0euZXAnuTMEVvR5YbwvC1EzmUpN6/mbIXBbvd9N6paO/Ooui/zHq
m8iEdcDrZAjnJN9N8g51QXv2hWz7UuZ6+vuYX87Eqpf5dC7KQybz57BXMWATn0Ca
TcWrEvVtnR6/GhTbEzDpGCVPpLzIqVFH8grUsVHlpLsZGkB9FHISHgJmmBjIQ01f
HjUg3vbNCq97U/Yu9jx8L/abPA/ugNV4H6dGriqM7WweoVzBIkfdcNZiIjbgXpl6
09AhUDBfzrkVH8iBsvAhTXtXbSqOx8BI0wpImb26dYBBhR+0NKy6/N3iz0QJWasF
kR9LRq4ff9zUCnRfhbataWWZTt+6NUW6Se/2J1+qFztrIIUXgZvon1DTH0pCxOja
9SilJ57AUwPETAkPmytzuRJAQnhtEQ4zJQU72cQ+qrOCh3ZPn8XKfBs++k1lhdD5
2gmniU4I5OBZtzOizFhI3oEcZgMXpKzvpbd4j0NBUGIRcYKE6hXfSIf/VjtsWLSD
X7+XQM8jt5uw/XLaDTjQ5XZ/iUv+9sTd6Mm9GA2vJteGx0AfBpkY09Gy2Xbon1NQ
qQE00jUUY6IIpS7XmdDYX/7L2gvSEqSXS+vXUmC0Pv4OQ/GmUOZ8g+0JloH+Dk7w
S+NJIgwDQTgSZSOIwwPWW360l7kiRk+MxsrPV0rZszIa1YyXFd1r7KyJnOaPsFfR
XOkAkOJlIbeevSfnkE85ngRN+vht1m3NRzG4jG2/GoRocLqsbmX5F37/Rs4Lc8w/
h90s41zAQK4XGhAzp9awJXMnthvmDSWxn18MQuHsauOS8y5MRALNFNlvOb/k4LMA
lxlRGDyi+rNHRz9UNoIXgBoo/ghKanSoO8ZaZq8Wcs8nK3ZSjBIlZQ6w5V5Q914O
KE6SzNCff4xHgSURciPeqiK+vHYrdxwSw53CRFGAu3+stHc9eZUetF/wT1YdE/d/
FE99rrJqyQ9VYRPn/wBUG5MPE/TwXE0YZeJ19NvvATO3N4StW4YcbMZDgmm0+geB
qJVWHowmkHD8Ncx/0vfSO20BD8B/s5QK4bUg+jZ4fzqy14F4mZNzdM4P5Eh5HYbp
hd4uNUBuUg0019sY0l8AzFDFFatj0RGCnE29nw+P3s7CBvU5+57FxGc4GvzMngBA
SVgRyDBj2ZD0V7VG1T72xxXAHYSvUXyGF/EiVcGvkLe4SD4jiZUkQvkvFdns6O2C
Urp0j17x1Q1vzwSWgeyDgbBtCFsK1+U12Z+QmwRL9QZ2NvzGlXJZitfLL6dr/ZBN
lkDkOqF8hPCoqbHb0Dhw2gKfxQ66nhb8YuQgDQ0bZyhcoe3XpQbDIsLt+8fCClvd
lo4lX/AW38pCDZY4ShhkgkmKxwh9cvgRL3D4bEdIolCFWS8Xk9fJjR79R4pzbUSl
Qm0Exg+pT04NZqR/45JJmGajFD/K9FFJKiPFHc1IXnKW76ry3+qY1R1D0zvFt6LI
ikXkbntlu82za5ZzHsbLkbFJiRHzh+uWZpYrhOTdr+panOd3cFNdvg19LZ90eEHa
ZZ7dkZlnDastKKcxrdugyB63Z88taJ2JERFqyGAyI6JFxZ+NYReo/Jx0x0I3LlcY
teKxJ3alZjcCAtbdfpYn75RJfn1UxUj7TYIRjBqyFTtYZpQDay1e3cKqAPccnQDE
J8MCZ2w063I/yduS0eHpj2yqXNaQECYxPCpKiYlGTkofc2sWX5d0fQYKwQx6P/5A
thONcYVFYofrv8OVEK6WUPENHnths4XL+uaV7SD4yGyVIfxbZ3zISi02c1K7nNwD
AGbSgu/ur7k4T/nrEuAvHAeNl6EMXBsbj7+bedwR8Kyd5DmChr6j7TPPm6HFG3E2
fthxzZuFR+HbNnV+TUgp0IOu2n9ZNZgcvKDAFqL9owvLsA4ic9xWOsYT4p9mLCKp
WGQCP9EWS2p+WRiXq7tqy0kD0zGMW/ESQCZl72Ji0WzShgAUPGIUY00KRJJ1VD8+
XKIWZIB5PLORmf0NJSPTswG92XxbRurkiU+WiKu+WnrkKO1xpB87vW3TmQ1GlHwq
9PGi/RDVaZG9kCm+VOHP6Z8mjYl4/+OkljhAoE79d0rxTngSL5EiyeaT9EGfOxh5
PpBN4sOl0Id29d28Jbfqgc+hF8uLgtGbcAxURud/WXoifsSC8JtTkAhd9S+CnFf/
oj/rY6ssna6R8yd3/eQqAC0Kw/VsFM/zqxh3y49hmgKUrA9zRq53Dx09qi5QhqaU
tCnFPOPS43V1NMqVTU53PouwS51f6LPrfGhZWY5ZhjKHbakR0xEWcBX0pizxfQhs
96R02mwG616z5MJQDDwWCpta75CbCkesk0TAJuJ27V83d/Ahmt+QIgHAzsaxX6V3
aRhdJryJnnJ9ZqU2JaK/X5SEgIw2vE56IfR2e3Q1kD/6mEcEXBjNK5Jy7J/Xyt21
pTNF+bNkRB0/sUmD7w2O3c7N6/6Pok4Ar0f8jbx6pEaae3/w7MAXhxuPPID19xqx
3KXweRs/mft9M1DurRbKKuTa7KATT9K9HA/8gJ/LQiJIqfvo7Nhwm0oTj6wNDxwu
eIAwHWKWlKd4SwsGkvkz+qHoVINIPyEw0a0g8t1qYCgAhPUzqzFRzLiff7Y61W6V
sjETs4BfC55SlN6tkCtA2L7zsjVsr/gIUj+gK2VTKPfs3g5o06hv20hqOp3iGbxN
OOplCmeakVEWnRLMEHgncnNnGy2CF6f5iznSZMquRYaVkFC/jBAOtj8L5ozmPjH9
cLXRcS6IrwdQKfy9vUaX2AIjZ8k4a7qZcW7mC24z1LcOH2rjb3xNc4VEL7iKNxXF
D/Hr3rf7fNFrVdBuYRtOEqY/Kc6aVJZngPUNflakWW1g1hXhErXkS4etYtFna6hq
+0AyYXzC0RR/qMTLI6nV62XrynN3FylKxwqntCdryj/SdCtgLFPKKC7FaT+KDL65
jy8xKfPn/uaQTkzspqescnJALjMt8zSZ2uh/mLMkItBCdq7zn0BtgQuVZSGA7n9y
6bT7Hm8VP1aCGuUdK2I4EdgBigEGgRk1t2vYA2IpxyYg0fOr7LxY+Zce8wBkLaOe
Q0luO+xxiTm1QmdqhD7uRgMcE2T0ivPcSURM6twFbA/W3zKWcULX3g3YZ176ZkRO
5T1u/3lLmHfk8nlfyuONs+K6Q6JvxFBOh+Pz+ckILpuxtbJqobHmjGAiRPEeVPlx
qirQ3k8QhX00t7HRYT4wEG0fetGkeZ3X/My6MEiZ9+SajZYw97CvsjB0OEySoki2
L/VRJWUaSu+6FxEBVQ/B9SawSFfJJCWmJ4JnHTv63WU2qxMjk3vj/AVLERe7hcNA
cEaoIf5/iiuroVundS8GzF5i2H4iQrc/+beteQtvuqWyUwCiWT8WGoEvuRWZeyj+
Gd0k9jHNclS/wxniF9ENt8xtkedrKhuB1emU/Lt9Q9pWg1zDOSWzrk/wcIqgEaGl
T3YTZ67ThicCyJU5Ent02hjnDyI6WailFo8LLzD+zRBsfFDU2eWZM/4Ga2UxHWEw
w+zDKAIaf/NzPSUAh9wk7P236CGhlqO+G0/F6tlWKZ0O1nY/Tu5T1+47q8hPAwyM
O23hnm06ys6Hkqg+yu+FE4tKAnHto8tvqF93T1HdNABv7RXp4Z1pwmntYQFWI1+P
ZQ+Lqs+e3ro3/lwqyhki/K1ACVw206mJ11dS7oNzjWFl/JWoKJ+UbCIma7/UDKdY
BXddCQQBDAZQwQfVmdHfr2Slo9Wbfwt3GZctyD7vwLBcrtjdNbE3H26FWPqshvAG
1qJ4w8QbQXbyde+C38xw+lEHPSbx5qB1fGmgg8VE8wEmeyvskwyomYJZO/3tGM0S
FW3Vtjh/s3Cgm6UnA1BhocriFw+mqkyU+N/W6RzjPqL2jEzYlwbRdmqDPXB0j9nO
2CJha4fkKKGsPPwwfTFfgH9acAKUAuyqMO918vB7Ao8R0/hQChgybieaTgb+4gtj
BLQFLGnodptjZsnX67VQA+FAHYC9GCzvKnUKYdchJ/N1+T4AdvP8qg5IIvShyrPT
NkI7uIOHF0/B/8A3pMTDduV/g8e326uQsxLWVlzLNC7bug5gzZD5QpaPlEGYV8vk
eINo3WJaGzxy9CbmQS4aLjTmq0kAMj65B6bWA0SbmQDe8ibmeI39q+MPAr1Gs1j2
AEuvneAP9FY88x2Epv2zmmgShzArT5hhnqC2h70fZ7eePnNtkiCICD9w93LEXFdq
2PMbbSXWuVg79Tx/6qeP1pObGa2W18Hjy/oawvl4kvQbcqHOy9rFDR/52QdPmKmO
jwDLA5X+e3b5dss1cIB/6B74JlsjJkVw/SELmIEQAtsopxoO2CjLUNyaYaKtNbjY
am5wTxtoXWy9w2jKKe5ixno75wCl8wEkLTn5dm88i7PWP+9q2WbfRqSFXTSigxxV
vKcUE5vRUaBgkc2+y5VEh5rPtrUH6GYlKZOIB1huzL2NO+VVLF7Su4hBVU3lpvhh
Kn+jz7ZzOeO84B3zrjqsqotfl+pT126+OZjML4aywazZ6s+avyfybC9Bvq+4dtd5
0pRpuhIe8voSwv0+L6eZ8HR19b8ifyfvav5q+E8FG/5ZmUgtTXE2XURIVaC1oVm/
NtLqWg1HCFrn7zrFkiFtf7DGDNFVuDTYKzGNaCtBJ2B9LAqs8KsWp2wQGko3H1hJ
fLrHnjLtylu37vzwiC+Dpw20Hywk7G8oyvE47MRdt+0SIvR/VPshIR6h7lYqwaz5
j8sjc5ujsBg7FoQNLZLXNcAD8M9PiP3FQt4Ew6Rgyaipq2qGk9LD+b49SOABCcn2
OwhoREy0zwsipyTifoAMESFHShFtFvR+Wup1IDxskngDvcEcmW1PQoJEXuuI2nbF
m9OPPserneYYLqShsS3K5XN/Q1o/5bQL8zrlb0JwcDJNkaeDMqHBMnjr7rzlAjyq
nBT/JmhreGkpwtwFC0KpbP/IHb2JJr320jPZVt+Ja4MytQOpClSXiYxGNL6cJLqp
wdSUauMV9UHqgWoW6ic3zMUXSk5ISUe1AvAv8VCabMXmDyI8A/YnGBxI6VUkJr1H
/m15rGDlebcOt2J3QyCoaPTm95UB47vTFWFyYUaIdJYrFfGr4BO1SrUGLv2GgL63
7vfZHf5bWku8QNFG+ZckE65xUhscsYziDKClyMeYBoEEfj259q3HOjXxloEejv7V
84c9tF+aFDT8vsDpvBAFDa3CWwVTb+D1LdVyu+qaTiDyWCyX4GXKCNwqOcMMR9Ao
Zql+hwDKaib+03uvG4uWB1bzd16hEeQzZC8DpiIXwQ19TZCB2hwho43hgdlbpoEx
0kKM+kzO4CRFk4RWAC3KojmsRWZAQ+4zMzbvXodrUWnM3CiWORrn58jFvxx4VUNF
5xps/ktN0yFCUovtTA6C8Cx+wsuZ5mPtjbZ+I/0VvSkfC6hh2Ui4pj8uGZpBetRA
xYl/6wtqHA8wbZZC84Dj3hjzEkDFnIUFqBqrUkTur9siEgYoRfx2Tg3TCX4jWu00
m5O226E61iC3IJlHS4Tk9+yxRXhHnukQseSmjskiCyqXYwmYgYNFLy4WVrXJjjIR
3YQGgPs8yf+8X+oSXPIjE6pNgkSCnhBWbePwbwMjMLCqpkewM2ttALZkP+6N6lhL
yfd8Pm6TsWIevoTwQZ5n+fBl4b7M4H0ZMAsZXbiUsKnxeD0+StcVEc8mtFN4C5Dr
KIyRCkcSC2M+OgMEceb2u0FzCpRr6nJ+M2xTgcbtCkrr/KErT+uEpJ9XJ6KMDUyh
5MUQxVlw5fcQORzSE8wXSsWlKZA4tfGu/jGsjzoTos5owrdMz0MGGigaEEGIeOa+
KpPPjITBF5zGL0DOkgni5+B18dSgIC9QKrASi4ufiswlrioonUruLwWLseDBIW+y
VG58fyDg1rDYT895sIVFNdWfmmB0PBj/129222cgsgbvvu67lGnY9XrTDJK6nGXJ
D5VCqlTcLhjblhrbvB3cIEriJBa0auBffNthvHOTl+xU6I0zlAIcwyxa8g4XMYzD
tNQRqgfpTE0r+9OeP5TRbgw9UNkT6osh/nrBApeOdnaaI4XxmYdTuXwDu1VbzPpc
YrN1LMS2DTbziGT7ztKfhBLWfM6M+alc9vu5o1KfpvL2QFWR5Oxj3as34S0CjhJA
Li8naPUCbNBhyURh3kM2nCVwMN3PLNo4fsM/LReANTVofGDXwvtDyHP/YX6P3Cci
+DjuJ1f6DUdoe+56v8crV1JpO1cV/SYsmrAhkEk0hlcPEFTCSNhSDTTXb0ks+8ST
/mwEx1szgFqqhRmzfCXtUrPQ4XFoA69MgXY7C9E0kPYcAHaEyxnohC5ZvU3Yn7G1
1QBM+BnTV/jRnyt8d8LBrHHkxAfjEbJk47SbVB1qt0yEEAZb/xGD8yqVudztZYtI
v7uekx/3JtbSYRlk4qHZycfUGlveb9J8PkfX8N++VxJtaYx3VARkQOjxRyVFRG6P
pxDvoF6uPeHMN+uYghcNNr8Hqh4mJiUZvBPRACW2mf3IB7ytsDwxbPqKDaokWUw7
c/yxrmDqaphQiHLV8QP2TCly1A6KuJBmIYnR+N9WVQQtCw6sBA4+l31JLMDLBzi3
PRTUxZExBcrL3JwRBRUkypy3c6syzqujQlImPeV1yI54oo2loBs9NZnFa9QxnLmF
kkhtHBt3HnrfpneatU6zaA9FoBrUCVp73GnTrKatwJn5/5q1s8Iq5VHCQkKHq+e4
0OG8dVXFQ4A1ZN49ayDNbDam5JnfhbgHoSXEYBb9UvsLADqBTjrI69ZB+uo0gp/H
I6ozsH/55jSVdRPihARZDQkhfynhhlprxxMjWMKgiSCAoNn9dMNPTbxud7pX28YE
ELXg19AJ8LcaJPo12SITmlkVFpevOtqmbLJNovjvrDwyqljz3X++jE/8kylzqg0r
DtDblSmpMu1rlFHiufgp/v14cWAYpvfJSksdjG3oy9r0yr7roth2Q0XYT7rB53Kk
yaRn5cEhV3nq8Wd2g7kdIBi09ylJi83CRkA2MlnpTM7nqmc3+O6ECVHvEd9MH2Br
Nw4SZDNfxXyG3n/K3ULWXkhmGG6ymc5uL3tqtFeFQRkhPwneucbylqumnsluUVhk
CjRMUzu+fAvOYUEpZ00AqyxdNe2Xp1+/KBliwhgkaSrOkWIP1c11zwOVJdXGqgx0
FcJEysze93xCIQXhq/d8ARrQSVgv20p1XuzwChyUceQeJ4h4gBqLmvEDYOni0FIq
EjgO1xAkiWPeqQ1vkJK8NO9FveT0AgMWAJLDxMJ+EkUoF39FJQO79ypZK2FiMmbE
K1QHEhr+mz0b7HGP68SxXt+qiF7KU5Uw+JmHi8FA8/+0mwXiBlDpL2CiOumockfr
7G+3E5VeSHVhLDtJPw04qkNdUPOOB+BiUExplkB9kr04doWv/Wd/NCsgbfQYulLr
AxMfCYTomuCAyCv+KGjCwgTP2MVO0CIdIWbJEU5fHdVOiRba37ARERGJ0KPfjo6K
YHhrxJ/HVML+jOpvaaY6PT5PqvRGDdzCtqL0MUzmwLrDvjLQzH8ZF9n+gGvtHFqZ
mxIaPc76Paq24i7DL3TVGksaKR1I5q8ORUUDbxWnoqbDLg156eImS6rTI+YwpbsW
4KXratBmn434X0CD6AjEL/yU7dEJA0J0LGg0Y5bnkRXgCam9PFTD00mAxT5c3TWM
MbOdSw4clw/zhtTbyg6lTZLCN0FnzGGz4oAj5bGQpGDdkzCeTGGd/uElGAl+Mgjq
kIiI5hfQU6h/ISwSzKv6VIoB5A1SUctl65l7LUnJnhMenZrAwGHh/b6+kCAPvf/z
5R7uieGMfYz3A4QQN7JNql3w2FfKj26quKgwkwr1R3MA5qPDm/c0MsRcWYchJ7Nw
JCWh3BrdYBDM/qc/Du7AbeBqwFuJBjiGgfNjl5ddXjDPnNSif5+WSEIrLJxMymMa
+fotg03pll1g5UK26TcfIyQturO0J1RhGf9RbYZdkiW3vp5VasmLbwrUVqeN7DmT
lCVVMl5wXWSTTRxozRa4WYwyhshiGShbK2+O5q2Yn67VvWNwKLMphCLTPTnr/4m7
IzNn6865VZscW+gcMNAQWjMrOWv1GAa155VUbAjyFvrVsXesChR4xGB99J0XfQS3
P7OcsMEcKW13k1K891lYypGeLC3X90L3q6xpSot4JtOBcZjwKRKy90qSc7hKeYLB
uB+1CbKMEmkFsQSU1dJGUXMUJY3CQGn/XXe5IuRyTG3f21iG1JWo6KmDsWHIEeiJ
SPhfPgWPvNMAoxr9tJ7Dq9wjhk1zA+A5iqZdUNXoMlXP4ZHT2S8yCrKjtYW15WdB
dcH0o16tNqY2T9Zkvnm2wamK6B24/rdIu8FQ0Sc1o/ayZq629FiCL+cjn69xGeNL
6LKPGCQ5808ci4ixK0MnMp2xS1i8o3nlvCfUAhaLX96Dey7SbU1L06u7csMHhuGA
/CozBmdrXH6kPhU+rYLwyTnKZjjrusijamScy2gsikBWK6/QDpKXFHeLHIrI9riG
ttt7TqKHk/k1hiSGv+fGNLK1i2qowRZRtUuPKrxJ+sDEFtk4wVqO5hAXfQ8Ll0ku
iBsN9XxOA9U1tkcozRtJYulys1yxdU+LgAyAVXcJNU53YJIH7cfOwqT9sT0xKEBP
LXJA0srfD0jJRm6/xNyoBzS/p5TK6vCAIFj973x17811w7wC4m8uvUiDC7P1ltgt
K9TbbZxI74i/1ZV1D7Rlt6YxU5DgHgOppr2zes9BpxAh+0bz/2CanyvyKN8Eq4Ay
z8fxI2AS3urplGWMoE0vHWh9IdgaYrcy0F014fgkglaI+LeKQ72LadUAXU5ajDos
4JRWZNDLWDgmFZIaeKcY8U3aRP1NmUUt1rMsEXHUEaWfXfN63YA/7UumdnhYh7RE
AUlBe8da8y5TKMRcvbsLayZkJkkbaJYRJgTCykFhqtfs31WPaevBhBD3/Td51NFJ
vUd3pY6kZ3PFVMgw6U4kKEhgmz/yamwCsPDxABESzkJsTX6IyDbiX4vY96WXCZZb
n/w4m31EqEL1Y7RRJgS8kCWaT5+Bs9LKkdjgjjUdPNiNIkNlrh0hbFU9xQV3eCng
WulY3rYMQu1LASHUtwVEuiXbe0PW0oAb5tVQsqcuTqcC6ZDT5rWEOHLVvXh0WNBF
vTc1hwJtPRGvKFceo83KMBWzIYEI6BnpYMWojnjDcDi75g0eS+e8jLs24CicUQu+
xjRO3V0fIXRU7ii1D3tSkEP7TyUPpjySfOH+i9q6J7+ZL/N0bSd68mlkOxElBiFW
pZFh50aNtxhj3IblpChWS8r9NMu+3XdKQORxRHEFVaH5vGYsiLekE2H+DJeY57/u
sTg737qMpMT/BTSnJBL+rrEB+gjk5dxmzOVuBAOpUUi9y9DLE+nZHzb4j6jUkzuT
8mMvyrUGMfDjf5l823uf7hadrKjSwiWMNC524LMi0SSrz2A5fOq8W/3LqqISZAx1
H2physTEZIhsULh8MZs5tz2V+TyCcjQXrPONe85o8LCL/Fh833tDFahxYCQUqZJL
FbQMTw/9YCI9PWE/VziFCCj+JSZsdsSn+K5gPS29UCt2xGL8uP2ioFEdUkmUEB21
aE6oEQap10/bXjwfjKU9lM4sBn0ZP56r4fQMseJPni+duVALiu61ZhZTvhmmray2
bRiCXSfkxnCfQuDWchiUaV9nl0pfdsO/4wOePJhplpO+i5sqGN+Jn3jmds8/7T0d
AlqryS31eJgXMOQOySsb4pCIdqMxmQiVL46LQ/nuf9Yst/gGi0p1zUBR5/zib0Ut
RGmTH64N76bQ6pMZdiAy/EnA5DhIOenrqMeOglU8+5/V5b3HJZ4adm7rl7atuSXT
NqSaolulPe8gNueWd/v/1/VOBTnJkIb0GHHKXlHmTFPmc5GH3pqGNVpg2oef4zFT
MwGnzWV6ndRjRzFwQe7JjVj+omTqh2kdLjEOMATVY+l9rS/MDthkb5RYrjFN73lE
P9U+IiuOW9lukTo3mE309ytWJuGD/C1OQBCFvUsxRzy4Z1RzQetT0ZiSasYnCo+f
bLijGodEfNhZgYgdhRc6xFKZgvTbXTTt6cLwB7lpMmaGc3l6rbfxGWyvHkvzSoJg
Vblv8zBi1mSZAcVa8d3IVepI+FkRZ1j/HzPrPtpcwPAnQFUru0uka5s7VrkleRnV
tIQmaPSP+mmN5XSPlPdn/WXI9bLoca2jt1BRGpbQ6kFJdf22TFvKLuvD6v4okq/t
1KppInfainWfv1R8ykiEEg/M+2Exb3dd/oaNie0lpYMZW/sqzR86mHo6cLfX5Cze
womb2Yb2jX+QnYWn8W7au+R806zWtIXjfA5ASTJlJIAbNAk9llBVSE2T3+9tY6d9
6P1qL54fhrWGo2xwG4tOczpMwF+sDlzxANx0InqonhOWLeIAYG4dTQATCc0y9LJF
YPHceTbqVnU7g9INfx+jbHjV5KrOVKOFCBbiTTg4OKlPVRp4ANUoAb/eQXK0/0B8
+pfpOOYd5e1sRfmA9xxgkSCZKc5T44zChhZn5HWJl/+DyCwkIEdKgFMj5VAYAsAt
6UOuq718VfsSo6sdiHpVBmzsnOcxFssU3xTGbhAWZdpNmEbOdxMpNyLoVf2S/z5C
olXQL1Ivs4ykb/7PgGEo5XfYq97cj+tks/z1lyydolrj87HzwVKjjOpbb9slCldF
dMa77Xe/cbmO+tvSHsIAS952lgyjyPwyWKe4WH0msBecQUKsooam9IBkS2mfyR55
Uu70UX99FoWn8hZTcYZaSnGtJ6rxH1ZbHJE7h3sy2NBUCr0ueei/6NTHIw6gQIDs
zUOb5B1cbGdHRnu0jUC3gCDejFrtPKJaij80OOvDso5qg/Du4ZRpPphC2Ie+THEb
GQZHJAxhTzGA6wq7iNmgbxx2aS3svZkDzmL9EsFTVvu3I/kP5/gr2++18Jf77Ll1
MstRJanxEBrhRZ3vN8EUKD4+Gb8orkSNEATk5CxPXT7kXVLSRyQmwpgwk9t9ypFt
KrbZJ3qOYBUe20aqAHvWAY6fGAYmkz1U3lUlUMxmS3EQPEI832fJ5kHZjgT85Te9
6YNQw7BswTlt5ppjhB0s+DZOyU7Jz4xerua8Pvvkz1gzwoRoLVdNaMJ85UPkhDb/
Ad7PSrg8RFD3aRjcDBWz8X3XYuenV1kzTo0lSclLlArF1qc59a4XaPTYx2P5lFiZ
J1GseIbyNbc0bIsElQWagTMus9/H5jPjnwphTyazSifc/EQzV7sgpEkYkqT114fX
2SGhzyI60Vep+d72LtBVp/3jxEQ3nJm3/xhkyMQ16EtooA2eEUW0GKaa/07kkecr
2Jj2GahVwKqQzZ4TBm0XmCm2Kz25BkYc/N8YDXxMX67HACNPBw1VCWq2S2OZ8CDA
SzO9gzdMtDNdVKzv9e4maJyQizefY5bpxNMzCR3KIImc0tBIuSCuo6t/6EMmo95P
vfXCO53ljiGdbUwIGtawClxfdVFzRgpLYR3+KKFS9ZfikMAFxyGV4TwBz4cS9NF3
nly1+wvTdYt200CkNguW9pfcT1WAC4fTv8XlbZw6fHXuv2+u46vjBqOZbSDqYxxB
IGTRcLTcQl8JJFnk9O5FplT3q7e/P6+m14I+2dM9EiqCmPt+pFzupxvrYKudtjQ5
snceu6u2zAQYGC/JGwybSGBiaJo9Y/9ww3Spg/Kis5DTPKmaEq07QvNRdPIznW3g
tM2w40cN8C3z/lkRDKWe9pm7Opi8cjyLAOOSvEqVCGXS8qp9ia5Fut/n/dJtsTPP
ceRLBJM9NGS/D4nI8AYG2jdtJX7kahe9JTyWZtm1D9zNZEyrsDJM3OB+e/kMY50A
r70n2GIlBNeRHZpoIxI93HNGPujv7NI2uj31sFeTt8uDMfj/BQCD4FVmHTs5hJ4S
np4XF/uhzel+W00kwnBRBsI9eUy4bbVl1mkG8ycQg6OdyQVk/0+CwSWZVb8H1Vk5
aYnTjUyZ0i263BtgV+IB+ijhaOavhaLQTlwvnYVoPcVwZ//3iivG67JntnUvyylw
OC++4OKZfwGGkERm7olwr8P8AtBzzXZxJSXphqs8qoTn4qHOe4shXmblNCUxF6JK
NZmKJF77CCR3mtp2m7zP9Ovz53dLK+RDuKFQfGIYdsaEci4uSYRe9VSjqUOTlGVf
Rud506/f9CRq5O3ezbdDSmqnFrxLfwcz27NmxvjowTkwD7KtNryCLHMG1Mo9ZjIA
GIaLYgIwsGAvYFykYUDOpF7C+113Zfl0aERX0+bagEh6J2RpX5LJ97Uj++OAhtQm
8gL4K7A7CM38Zm69NtSdeH2q5LzXn+EHbhjePrV9GYLzVgjXFqZla56Ffy5xjieT
6oySHIrX5dgCuDC6z8DHOoWzM2IcN/J2G56IkZjqK0ZuSGuFX26xsIqDWH2z+Yh2
xKUBPd2/pk8YfGz26vcIMFKHARj2Xynn4gNjqWT9S7MhhGEIJ8MV6NwYIO3GtvFw
PwPm4diwT1jebmndsAy9BT8UmNEI2Q+nrjs7Vgzr9K0XT9yILUUkg8YnDnjgkN7V
wiSSPOJ4tVuNBvYMwssInr0uxOVwFH64Fm6wsrzaKTvgROwawbDJfyfj5OrRGcg4
OAsQh0t9KkkGiUGmuJXljgtyBoLCWGgs1mWsFnBUIIMhpst16VL3Osm23pu4FN4T
HC6u0GLKM3QBfRJ0+wDX86A09Fh3LHCmeiyPYNP1hTQ5AXYZAH7USbGdgWZdCRkS
p03TNUKA3mejHI0+Do1Eqm295D2+WDjj++AFe5LekME2SxcLTeiz4xgqpuu+K1Wg
yvTRy0tZmR91jcyDOniiYNBPlfNJqGIPGjjDUMQzjpANptdk3Nqg9AeDkurWBIJl
KC9YX//ZHVcVHaPWEUCHjv6FEKtjKp5Tl4MoofzB9o+jMi9bFJAFt136hKLvlAmS
cLZjk9MHA1qg2o8Fy91lM+bQLZSo/PE4H5dfGL5ZG/ISSAJM1ag6aK+J+1C0YdhG
0IDyGqw/zaQsn+Ma1Hn2Yyc/NBXVBBkuPzXGtrTPn2vZWFk6dPC1JcJzqlsiiISb
Mkwu5bsQWOuu+jf7reQsyBXcCCN/+O1JKwNpgalUQb++fJQXKaoG1jlt9fSDEwRo
WxnfRkJUa0Sdx5Qto3KLP3av8rCqps82lWkXu8SX7mxQEXEQcNo/d4zBhn24hZRH
HPJlFg829ibuJ1l9f+yH3/USTbOyF/5AgXcOR3tL1N+y9BhsEDZKr7V1ev0IDoue
p/bDrfDu7+q2pOqY2kBnZ4gQKICEM9Bg+Os4TP9izsWRkmUK85/7tX/7feHxuLhy
ox4nX18ahvl20uxgCl/HyrgiTEEqNohCnM68RoSWGUQ8WdL275wIDk0Y7YKkE42D
pnOK0Bjmxp81Yvs+icvBBRnh9FMZ4eTgGIYQy8KE9T77W8FuJzmAOwju0cfaXmBq
Q06Nn+ijuxcC6Uu+eHIuy3nzjRCa0YK8Qq2XlKBK0ldo0e5Bv06Y5ZHAf0AmKAeY
kQtMEZoc82B3fkc/dJIyM+sHqqx6PVYS/EC4PtlT0pCO7HzflpdV3zclKz4IPgtj
/ayQFzj+qrC1CyiaXFEbXLvKIy/aixCwGhmyYb+bXepa3Wil02iMxx7SlAciL7Ob
b5GZqVMsu4kHuxcMSeVllqff0/1km3u+XuwMjXgu9+bRKggKg0Km/XRltkA/bUDX
Dyeb7AciaidwEvLuwzQzvwkfQdmg9vq0erm/+rLcd1BKDECABaO6AAzLcT+v226y
5Tr+CHjdNnzd770yTzYIVebYTMubS4NdPkuzpMrHJcJJvuEDAeud41UzQ4ZcTv9d
TdIwSe0PfkEjeeEB3mDkXCyeFhxjoCTpC0SVFoSSx1hL55mm0/uoxH7d8ccYKyKA
hKr5X1CdeMvr4DsfKC6xMnWHV5jf+6VtwxzG0HPF17tI3W5awDTNUChBlddVRNiQ
ITbc5LOouv/5DvGbltNkVG+FcK2rCvz9bEX20OcwcJMJsJR5mQ5OJ5HNYPPjlc85
Cym6QYDiGCjwg9TOvhhjyTTTb7cBJQjKu9lskITW/Hl515nEgNMMvyJayLBB15bl
XxKNfqTmyLAZwI1ZWQVLChtHB1W8x0UA4cWPwiHjpo8vBXnPYt34nvnSjufi2qNz
BXnK7nHY69+0rJtXiMy81KEDEqnNt3Cy3RtzITSk/ve6tGqiRbWuQpIbNAo3a+MH
L6Nhd51BmJHTLAS5mFeoDgm/9DTRUxLRH8gpz9Q8Ify/nGwQE3JnWEj9o1s6aok3
8X23df64inZwZXb0iZLtM8NwEPEGNtqGeza6mjBU05qLxdsy2KFB8sadTshnDMtT
0Mi3+Qu9uBNSmxIGttgmbTLqhqxTMscu6JMAhCH7GY2Hy+e7UVQVs28GG1T7pfFK
cxJcgOCki1T7nV/y4gkLYmoyzs17lUHw7ATR8mceUzU93mMpdQHAPE64vAYuoPGI
Gg6rGpA7FALC4GK/hV2sRR6g2j//TOm7TG9T6aVEV9qbQWFxllixb0eIyXuSsFSj
PvmJquRmfWW8gSWyJTYWsuP9zqOdP+gaMWKVHrM9B2XDrov9iY1Efk4Z61xx4ayx
QA4vWTZ9Anm9yeppns7Ef5DYnFprhEwga0HNxIqYBhc9P5Gc6bpoYugJZl+monZt
VqZY7KfHu6H85GEbrSKF6QFPR72Q/I3jR4NRa8gFnaHYNHV4r9XSwr1oqt5nzhSQ
k++FDFfb0BZ4R/NYUy356m6LRcqM2ENpXj/rMym/RTATukiHo++aOKjLRSqY6WrV
WA10GrlUHMfKJwjA64qbmCPh7SQehxD4+M50XHiGb4Hcre4r0vCe/s2DeAabz5Eu
ysJpbWPBaifb7+msapJCwVO9JNmswwvXQMLgTI/3G/qhPiNoD7jzJ9Rkga/KTfIj
3ik4oX7WthFEA4tXUzDH0mNaJwcjR7g7tGCfH5XKhgtqAW5/KsIit9iKHmBj5pOQ
pTZjk7JLGrCpJNd0jyb1pbgEHzMxeyVIPvjd8cjDiPZ2heOLEu5aYzsaxRtJ9j2G
uLtkDJBIKW+3IkqXcz2VnTDOi1DB9hZWiBNctkwo2c7DWaLKWhlTEak1LyXRk5n9
ZE1+I44XuSslxSh53Sv92rn2mek/NiLsKH4Lse+OR/3zytoeO6TNUm1JfoaQVcl5
3RPqb4V6xSElQHQNuO5B7ntNWzpTySxEwBa26J9aDQ2cgn6alcvenSIFRIhqRN+C
8nC+e5Vy1d01+w8SDPRhyr/loIHP9ZYAOcQiJrXycj3EczOMy4bNSlhh1d0Dsqy6
PhxHiGHMOM2KSDW2jy3mpTVl7p6mEZSQIR7AYtoP4jlRxg5qLPUJWtN53t4VRGtg
Fp8wFokzQuwDXvif7pg//kQn3J+UO30zduLm2sACHTzlOBj0moWicJXx/6hWu2z2
JoMqNEN0H9jgJWkhOt4o5XbDu9gz+cxxpq+tELmsRxN6PPmxYf/XDa7vPZqo2Dw4
mihVULMmLHC3FjCiBSH5ou6pT1lCS5SuX3Nh+ZEpWCNBR8EwJ3VSaUa4C7XnS/f2
tTSQlqnebSzZVcddV84Ha0gDSqtrM3g1TY+xtggsSBxflVeVpumKIdBABVfE2lKG
oNbYRAmB7W574a0jKUP+7dpvc69h8sYhq1+RyWJlk/qIPVgPX+tg4OpQG7eZXi14
/NFfXBLCZMWDz0PrucKP/x3Zg4CX/+JJJ/f895ICKk/f3vZ71NVsNMZccuyC4TKA
q74OWXgljZUqLEfLeiaDUAb6zUQk44ObJsTm3z22tCws0FJHMNeB0q6lTOeYcZiw
akFAobvMdrz7I5HjTqz2wwzvkWwZDMoiqdnpsXPTTK/oOdqtx2B3HDYTQA1n4CDZ
0wRWP/Aa2jjd/ZDu6Kx8vD44eLwgGlM1anWevndWf2b9JHTbcsqErlxp5PwF8ed/
juc5tkMXOqS98cfmomgDBOLLNFmeVZ9/B0S9n2730C/EmyH5y0Nh0L88Bupcc2S9
vo9gTlw4GbjfOhwQJZmcnMppQPH68gqGh3s9AU2YZGUTn0IOcB1EZMbb3/kgeFWP
qGFHa2mCxSOmL5uDx+LAWghDtinTN9XcB/p04CS/D+qa4wMKpFNd0Y6sKS9fn0bU
mfk76ifOPhCcg6ZonNl1qr1/NTAkmUtShBhKkb8r7329b6cBRNDrFhjZeYNIwe3r
j6j/jD/+4ccqzjPZ94uuL7oIri5z2bpeL+h8+DNjXuM3EBxihMwSmkbYGiv8GPWK
aYShtA++JT+JMqFUDJv4B9y37zc18n8LCd+6tuV4k+3NQaeTfFX17IxRhLFedHO2
WW7hWI/J9+5cxxKuIHD5FHe4uoutFTVn3V0BFuSj1It3kGJqt2BqE4KUiGtnhBaE
DEUcWNzRif6kk9liwBLpdeQF31pJNLvKTVF42eCFTECFC8jetdy471FnfGMOD4hu
MocNGl5ynZAJms+9AKO2PTdtFlnYSVE6d2TAjPvTdlJENrYEGvtjFCOTIXdU7xoL
KywmiRQpgiF/d2SxnIwz5zO/w8vQyjrDRUurZ14kScyaf/5xPpcABQpE4+H3EHxI
sM+70blHjp1Qv59PVNf9DSZidWxMA1fHLdPYRaifAhlMZzz2IBwO77I01aPXLJpE
qaf0I1kR+H8mXT3TNN10AIDT7fckDM0kmy8PKoK6b7Juw6lBw1Dvd6sUc4xmZ/69
pitocqBl66zPkzen15CPntv3rhv18R41/UStHhjJjJ/IRgG1bvqkJDdKV+GWZvR3
22LJMJuP180wxm9imvMUmU+jsSYmFS9OoBWapbjg4jQ8+rubpGs/8YbyIPyD5K0q
s3ZlmCrPgHbpBjF3Ni574qLG+1A2ngTAVrjQVws5Ym+Pxu0gYuCBGH4KBpKvdOcp
apbI/hK9NFKSqygGwvOi+HVoTohjnhw4RdDlteR5zqqN5yLmzdqYAt87K/WNHajh
BCIAM35XNxKoZ7+1j7Be2pBb28pElf/9693Ry1lFRpRyOyBwfHm4EPpF6nFuSMEa
sYBq+R9OaeaIN5VSrkt1YLwgtL/u3doq2/gdnEO7pIIM3tRj7w5hqRQRg4dvXg3N
uMLigsz+Lr0yryMI8DgZjyMNm5WfuYmctLtDYt4WwRp7LXFOQI6S5RioWHpgyJAD
EyeiIygVsC+eZ7ninUbOzAmyan5dsUOgR2dYIh1V79XxmKahVmpgL20n4J9p+3nw
9Pzl7u8VCvjxeJSv2RE43bj0msMmkSGaYTZbkExkFx/J01shK4/HciQJZCq6S3sb
XuyDFxK0lKfQ3jbYX/lmzJNcHGwlHb8FHCikfV7sKauRN4QwX0/YQfsQjiGVZSF+
xMISCFvf8YGvPRrin4xKjcjxN2JC/2tmBUXraPnIdcqXcxcVfPiF7ST/JO9St6aU
HxhGyKrAIHHB0c8/gzsbzBJwAGy/nbk/s+x/OcnqyCgHWH/DqthmueU5hC1yQbtQ
0nSg0WQ68Y8LnFZvOwrahrh0HzXlpSVfogkEaFXEMRo8IdfsSHf5xGkBdyXMB/BA
jNBqPVYbZDduU05qere5/TG0hweNrHRr8nvKQbNEf0FH7173+v3sQ4fUehtmo3hm
WjvO91Qqx1V3A4mqtE8sdwabTNXtfYcSm1G+6WkJHgJwNkJvPkZ77hV14syzJ+v+
Md/skojLkWNBPPbeehIyOp7w78rW5DMbgFUXmipaKLyEweGSm1So29ZB+zobioM/
f5lp8mi4oYw3wL0xSu1UTmRthlu37N7s6MJ5mjVjQCq2PS1uFhNQF/Nk+g90v42j
x+Bo2PQph9/Qb+e/w4WIyZwhG+YD5FH962EiAFUXGzRxFCMugcjBdp8uQXgKz79+
L+TE6Tt4sZjeviuy6HJILIaUyXx6F3ehHzCW1YEK/QTxQsf2ZApBcqIOSqykGrzd
Gs25I9Wl6kEHDlh4xqc4xwkEnY92MaQExuiN89vMbjvN/SBbFOMcNlmJIUwVPvz9
KADcxPckG2CdvHXkxcjwdxZujsM4jbo3xxK0Zhwy9g7GYHqc4/rNh4q7Npmwr/A4
I48WlzSYtP3CbMvFERX6b5LY75v9ZoXECmXULqA4JRC9CsD20dzfuaWmXuZcdJOX
Ou5oST6K2GqVY4vHiKU+dBzHGHbE2yn+vervpjqSg8/OG7uKL+bZWiIJ7GAewfyL
lPhqx0gFH6KJHugr68QiW9altXcpuDXVvnSdgdw9zaoHaubTlAHpc6YXuhFrRcDF
k3jbgNDGM+KpoDZIJfz6i6R2iaurA32jv2Wx7wWZxxQcDWtbcdjT81tQ5Kl5DyCY
/Waq3Ke92BKpQLBhVNR3mtP2CBCm5hKcxhKHQQHkcJ10x7b+sIV1i1DO0IqTyZCd
cuR8Pc7e1QFhlYxnYGodDZQaRGdcmygwrElAgZqLzhtJ/c1QcH9yVaUVQbXvocqg
/stkaVIOaFkXjGWI5vgwjQPaUw2mcGIhakhYzHxWGHrPJZWPfcz9D79RBGvsW9fu
N0ub3vdFYP/EQ2f9J/LocenILg2SDMR8iT4JnC1MY1msnXnYaDvrR/IVldBtiy+T
kv7WbKUSjbCX2yalbY0SFSX+zjU/fpcpIAn7Bk50puoraKACw8uf32X2OTF+/WVs
nKpi0UOz1nAADCH/0Y8xdZRqu6yuePsCB/W70WIR3qvH8BLYGag0xfASDFjK7WfP
KaSH2m0TRSFJ6jUmrE5W5tFJqrVxghmTL4ZPu2pO8sPhT1zUUx15vM9j8ZZAUWU0
3W03uRS/e6A6ChN77sTkT9WD4qBqa6yjWsDM9TqT9krPipOAVU88GSqhrfaNJVip
D6OZTuaFMdiIx37li7NxO3HI2pwjNjxD5MXXgDR4p34MTFu3yw+k7Ol5JjrRlbh6
f6gCJ6tceOSJfJ2JE/EfIwljTVOQZ4oGL8HMyuytufXOPoVX8+9NZQNh7jQIe7pH
awTMbhDxfFa9Vs5tLVSSwoYNj2+hdvqAx2eCyRnDbKADKsSesuBTEE4PMtNmN7Jt
74PNpS0qTGQNr7QShyVSGDgexrXS5fKmL8ahOyi7AFMLQZRQcAdGkjHxp2kEWpkG
YGys0rsuLlmhkS0G3ZcUQsBPfb/AXOxC/vvLgSwlkPlSpoEUVzjp22vx2HCEUrbU
ghD52pGEZuSPBLs1G/QGoLL2NOVFVmQqqFe31TIVLhwvbwjRJ5NYuBzsqFjSp9AK
/SlPbtEykLN8wSKUHiHdrKLvbEw0Y525AFh8iTwPZ6GLdJv0xTCmVGDftjA2RJyd
w7Vxd6F5iI+iHjTP3a0LwtfMr3prnJ/NucFS+fsNIYtyjfUH4bejKcsEcbYEcM3L
BRRyXIe8vO2Lkj6Eje/t/FDT8QYC2RlqeRxEnIdTd5/3m3MDoCM5jR55Zth+JhC4
asHzYPIPh9mEf5miWJ0k6doWO3j/Faia56/9HzN+PtMvDUyMg4iaX33gV4W2yV80
htq+KzZkQfOnXZo6VVhvHXiYNWWlyP2OrhFAREmjenWKH5Iw7bgIAwd63+jF5Okn
cES71orp58a64x9svGvBrwoI7+YP2znY6QJcf6oMbroMZKKGWhV5c++ywQDNyLQa
fSAbiD1QxXBXRgNJ96NH0UPP+r832A4UnIt1ktKVu/WSBrAMjRO4XZcM8y4jRKTH
BGATrotY7a/p80NIzXV8GpMc5m1+EQGUvYbUWvSakUaw4XxQrQhrwYE0lhJvWl0q
6qd12OJHa6gle0lcP8AARIGtAe+bsWQU9OYFFEYK6lzXL0K30dyfoOr5bR5G3ttf
lER5T/9Vw8v9PCkBE7Jlav49rbaVNXxrHioDEFYyPPZ8A6L45+D+WzU65A8PZwJq
Z+48wk/V7RIshJ2SPDF0zEhTVy5V0GOLDHyATQ/SsWCyWLDvAHfwGFAvqyz2yT9K
afvmmSi2eICor9Lwj78PR/WQt8lWldGqkLTljIp8ebmHuZicpBLrPVIQkYxMRt44
5UFRwDzf2Q4Cso8LtZSpcQg8WRvc6+mJhdv+bRcg8oDPQ2/Hzq9Kz84xM2wGFNda
Gyw085B8w3lvVhR8J/O/2ZPntGJBxplF0GaFSxwuxiNRdCiZ4mJlF0QUa9EL7RXT
J3qyXVgE9AlAu8SpJ5VPK3oWqfTBREEyH34yTmpcmG/3wvXMXkU2JUc43DpVMLta
l6ZsRsuQiQqJK7EfBVvuunOOEwjnEBgwZ5nV59YNko3rred39VNEE/g4lGZEQBTd
Aqaoie1zTuBjVdtPIMjJhBSyqHf5uSN3OE2stmBQGLUPPGE6EE0m9GrHrgdGFD5a
GLdv/r3WZIx5Un9jkG1EihhuwFRU+9udpaLMiiGutl7zjiAT3qZ5ZK4wsXnmox0F
X9GLZPWHOvRofMQ7znEraesC8uug780lOnIjIlSu3n2gzLhhbEsEYodeBO7/swRy
IBYLLd6omrTnLOSM7Z+w/nlSHAcFoGS9bPtxtPkx4SwWpaqp9E2skYtETcUHu6Ho
ocpgfpAE+3ryX25L/csw5HLZxt3O+N0/yi3hfr8/L3j7xqwOCcxtKWTu+bngtNQa
X2B+dbccK5qdM7KIIN7E/WYAxLIRH69OjqLoZrlOpSPjySFRLEHdE6CFuE9w31rM
fDbYhPYN+rghbW1yOADOmBjqvWFtw8iGsnlLQtAIXsT8dPj0jEVnjvXZD5Ef1R+G
kDOGeRxjB5SquBZ0/nQQlbTaOhj69xltMXR08Qpc8yO7ye/QQBBy+FmaX5WEmzxD
ypVtEnAYTtCOw9AgSy2toCuhyHpV+eezwa1FIxXocaQNR3SPCDkWAlHLP/pIqeTi
iP/zAKZME57BYtRdAhVlGxcOcnFpnTOocVorRoNIsYybz234owcoXGggX936/VPR
B2XaA9gOSu5fc7/4f05XhvVhJiZWozjA4hyP6Vx1j/y0feH3uYqIsu7EkufEqCea
AfR97ipeH7NAGCwkBdOztFkUqDjWeO5n96GZEwT1WCesQu2mhCR5nSLt1zS9yjMq
Q3TFQ77ySKZVbvfhryanwhDV8BDkVWBhPW2jTvcehBE/6hHjUebrdOjtSQJ77Dz7
7uJNskKVoSejgf00cMLd8TFC38gDcR+IsCNezQymJ27PD3uoeIFOMpdc77ykGZ9T
M60YFUSQrrITg//K0bmYw2WyueEpggxI+m+3htdVut1vi1cSScYOdN1RtCK/cKHs
FMvJwso2Er06C9MAtyyBkfRI2YHQtMlIgsp1Hqdvf/7465zXqwSMzR0lncW60mny
gZzreNXpfsVMBVTO9aEw5Lk3AEuWLqqHCl2KvKJSFOKwGuYiT+QDyknGH2PgxCy2
VQPM9XJPSNrQSY3JEZZ3wcFyTxYQkDBCq9vJEgUeV1wxu8MyyyfHTKbm49H+Ot/F
6HJ4ROT9VcX22RiOL6dgm4xm0gZ5HgthrXt9mWxDxflPZf2z0KKw2QL1sZt+0X+w
b//ru+sKVYFlb4xfVIZEAChbi0fouXWmtzefN95TDtcrjutLUH3a5S9+C+R7/HVS
vnVo8BpmqQ/OLKuMnAH7pRZfyYkxGoROuKWb95XW0JEsM+Kb1aX2Betly2eUoKmm
YtQ2KLaVNsSXe9JIrc65t+DuEUKF6+Teb9G/w6leAmqagfZSw4KBmh+IFXMRFUvl
fyOq6ZSRc4XZoB3nbDvO8A3qTFy3hpsywTjAeQhyHtX+e4iuT/jAU550QSBfqIR+
xhNl9odnwh1mFcMVlLAjPDdj32SwnmD2tLkD+0VXK8oU2wjxStxtmPRg2bF1uR0d
7Hk+37KMqd7KX5+IF1VBOEjV6W6a/Sp09ht7gZQJcsR7Ay82l3Day+dwh1b+77Ze
W6ak784bqH7+U9h4Ao5DblHp/f9wxTQ5+T7tWi14TmTGeQeWa3ePeKs3bF6KDYz/
2DSGCUBpR9D7Bhsqm8Gk6gd9OGag5f9tXVf/eipaNyYLKagofxgxBdeIHmMRB31v
fEhCzMsFkpJwUJmUVCP3LArdiq5MHYK/Qwlc3Nz9Yx9xkvudSQC17SlPsA4xX1IT
dYXT367rnsN7PHBm4sgQYUjiDrg4iPr9mNKnu42rjxLwv0MtpLwqG7j/u8wi0dOt
2V9CP4f9pG+TIyf6lKO3hNs7pw2mVre8bUIFZWntvm1rfAjWN9QiL9eV4EXKImTM
7dDzhNc1a59jmfpBqZQE64Ow0PjGVd5cv8Gs6e7Rr14+m0VMjBGvx2FLzXDqzxBA
+tAyC8UZyDxnj/mv8e6DqXCJoBjFhZ2z2In1m/M9gq8f9jNl9I275su7svc/qUwl
S1wzQbr46y2kREoLb9GUzDUzrz4jP2ynN/o2gGSKmIWn5TshLuy8tI8xr2Lg8NCm
cWDIuNziy/84XhdLlytkND+R5n5OrkZH86ufTVPF+HfywLSP5P1yd6YdlUt0Zntr
tX2QKpOOKmbnC3kIe0kjPbNNXwIX61CrleYHW/4GXvHjmRmSNUQAeRScw+DKT3dN
2PPiY2iaSPnuLP3nLUPSIXP7fgafWa3MbpnjC6LA3gXJ5jxfM72+HujAgfZGbWPV
jOhKNuy7DAc8QKp6b8CEpvumdy/ngnV4V3Poubt8tbEOKveEMowlVNH6STPQbTXe
2umE8NVWrDI4aVjjzDjLL6ATwrnWZlprE5wMKHcSfj17pD9khvFSdWlk/nsP4YSz
u99n4b1hU9eYqZ/ShX0Fx7VgOehPT+b7T/X8+L+pLHwG9MhV0uesrcgwlQTHTuCx
f5rgfvcZjl+bk8OHVzf38B8e4A+YtLtgeAA1hl+KlNGpXfmsCpUt49K/lWIUtPVC
XNBausAhpQqvaAgLHlvVBic5P9/9wh3WDOOA5zNSDU9GBF3mVikxRgyDkWM55EzT
ur04Ne5Zu4Qhsigj89yFBKQ8+AwLVmL/bHwm/3M60cFnds742DVhRacgzKtqoVv0
qb7LgqjGKFZbZ5n95KqSYrPq/30862tZqH9xSyJpQ8soCx7HfzQr8cerWKQBpayn
SXvs48gjrmL4VXu1NbKcLAuqW1s+WGi3OJSexEUoHbn4kJkLO2PJlHmNtM49frbd
lDZVebd6tFFsUqLH/3Amk9yn2qir9pzk+J3zeJ98RnvS2IKm/BPa9z/aLGiignXX
MutQo1512HKxTjNllHlWuwsDm5B9JFF7KDlfBQ8+U2LgTH2WYjFKDz85wsIYD/nq
2sE0j3h0PiCzFOeTxCOvcOzNgIbshaF58Mi8N7ZI6UwW+Yd3EzOT3VoygQH5WFQW
2TzodbAtqSoWZFarubc4FSto4J2qk8061fQDfK+KkCyWTHW4CdavmTfBwTgCMMRa
25V6kwVVTXOdTNEow6ArzyCN2WJYbq1NEdsAnPkpcFndQkjYkkKYaDB8RLSGhYgJ
i9m+VR7NblwpS99Rwi5sZ3wkt0WLeG2+p5oeHRvUVQZBUzGQxoYUKNAjI3jA4B/8
jdSqTZNG71lN0tSV/QoKrqttGl+mvbRaTA//4H3MLqDfrXXYh3SiZ1QdKXdpcm1Q
vKyVXcMUQJ+PKqCxAbZX2V1qL8Ln9pz/F0IEKsBlt/jYaiZV6Brn1cedzIbQtWwi
SAzdBdsvusoK+SmlC0nLIXgdjEYbTqgpRfcgvXptakGMBMDfqShuealxD2lzHEc1
tfhNSVM/mTzlWhPWai9K8SvVoZwAL8+fVgdTpIeIfpUb9cK+aKzCPpj6yqZjv9dg
KA1LzV8rvbM0mgHcP0aJRrc6JnckFh5QIyPn1nrFXSEMx/Lu3ULRJYfms6O6ponK
tMIcH29u9Rl4bxTfDjJ/BTXkyTaNWIE0qcUmCI3NXr6muZlkuOp3VPcZbtNlYDY9
V22brT2OG/BxaeMXEXl7KvKwbE+mHarEPlxHLHxpNss+7n8Hj5b5pb+zBQhzenM7
amFtQ0xz+oDCH2+bcg6xg85EFMriOdCii6JFZsXg6l7dZuTYIvWY7wyE9VT5edBd
Id1YipMYbt4Y03tKyUN6GdEJNxTG6+FhWsyXroixp8I6yugNM9rP0Vwhjp/7rzui
S1I9bF8tA3+RJlgGEG6zMI5/zb5BsnxKtuHb13T4jH3iYy+vqN/Y+h9pM5J7YDla
/nggN3R27O2Emu6VBMW2NUt1isXWFhu9JrVUfFciJHQDe1GMVY/9Pzxcb3C51p6W
UHtwW3CgP+9FkzdehhmZo9dc6RmukQ6RhOwatGOIYvff+h58DBq5WHrTZiFwEL7z
MRwFVgTWqWMwMJaptUeL7oVtDkojynttF25WQLK9yBfggmOU2w78RuuqpcEq7ACE
O5Tt2bV1lVwOmJ2HeZqkg1Mzw621296Gm4jhIGCPdG/42Y62bsavxL4mVkGDgmEB
eMNJnyPUNOE2c6cp42Jk0GGWHoC+b4a/p6Wo7fyLaPX7DhtvyH+66hkhkbwxE6Lk
SVDzIB63rmO6dMBVMNxWgQdjzx7OCxoU8RBToHXIoX/DAVd5Qf3rQ5H/4fKmvW0H
lP5hnSVuibZ4vXi2wKuqqmde9Zs+00ihc6vUn6C+ZQIfqhmZ083GhqKa6aSW+lX6
3H2OkdtTLKCjRPUycK5hZJA07QeIVh1K0+TH1nsCHAFr7rT2QliwvUcsSC3bvVSf
5n9UYUWBNz0a70waNcy1oamB5nX6muND1CELP4pWOz1oewrHum1mTwMZ8A5YlP1R
SCxUUwYBTvQcJxv3elR7l7HT+v/EXEAqekQIP99ja0Yzu1qKEWiBEiVmvNs759TA
AKEKPlyNljmA0gCLe0+K2SzPV9jjPJ9Lc8SOyWhcxuPD2HnNL+u2hSbo3mE22hpg
YtyIxyqki+h+5SEDboWbQ13qsw8IOZ3bcCaFCgwQk6rMKbCcN3sQTHtv7mIeW7Kr
uBO5k1XJ+gJ0/34xVdgBXzHfvBuc1qIzU8bLP7yq19da3TUwfbPhsPM9NM3unTLE
DjTMzX5ddL5piD8AzIYChyD897P04tW4QjOPiOxER9Ite5J5Pffid4NuJK9sGDlX
zUBoCkq/3RbJlWr/QmhCtskpHbOUAa5H1qwNBE2wN/NGGB3IBWw5PZ2c3d5776lB
iM84xQhcCiIcPfogG270247r3Rf0/ywFms9Bvw2GDpMZmIjpeVNLTyrvVadWC/Hk
iUX27v7HxQmyEeJICNaxdRq/XSUZBIli20+lxUZCeChU12kQKhjUtuhNBuC7FGz9
8k2B/wB/7f23HStGw3q+5QDNgdqDL5lQRFbSn6/LlHbEBEkgYRHVjVzHPtNfm+/d
4n5s9e/Ufh8Se8KCA9ixmKN3+I15dhKPBN6t5pbqsLJQe1bgSrpKckfqP9A8wSFD
oIfNyacsXg6jlT6rV5V7ldobgMCs9mr/UzNt4Lmp1z1ma+vGb1oC08KRxas2z/9Q
3vOM5G/1/VornmpZtIZlLsgi1jf4OK6qXKo8CscmWm5NO0iVjJ4W6QhZsavpfeSh
+qWKe1ntBMXAwogPNXV1Aiiw4BVgotDB/gMzNbSBzlaV5bgveABmzcU7RudkEQni
epcrIbJSzjgOuxArL/igpiZ53en8tf7eLCrIB18vHc8d6CgSsx6DYhcBgsePjGpt
sYY0YA+nKZ+K9pCoAD0wxtWVRUrA+jGEKI35ggVc05JmiGYWfECIDRVuQr7vUMR2
IDYpEMZRbk2rANPXdTIx5kOaOy4cYmNqsRzg0SmdZk7v315qT4FRdV7Lck9TQ2Co
hHuR9e8A9wrOAYE/FIc1uk1VUqtQUOnSOMcJByFWLB+8FKtkOYvPxFdRMgIZzBFl
1U7Jj1sSwhqf0Dy86uxfcrlZdGIgYgIlaUECDqqZdgLIsTVHWV8WgUVWrgBWjyFX
rzpWRhkGe/FuNGmhSKdOPOqkG8ONLw25oVa3/7WNIM322Zw4mVN5D7Gsk3/HtXN2
igEHrafX+ybrg/RIxIskH8OFQdFOwtGE2OKqoxm28fKRk29TtUL53MSKQE5MgeKM
Grf+m8JG9YBOSftRuYX+CsHgjHSuRryNfBhIGZLC0crKCjxmylA4h/PM01cxdVrg
YzrnRsUTNWS3HBFPVZUDkUwACbLcnPjlg/MhoeTckq+Na5zgFsShdAnBoAhVr7kg
CMmgIz1Y+ZL9eeMn6PM0jv2h4p/83iAL2gMkc+V6NIlumReeCU3AtQCI+6Nk3SLX
Jdj8/PVmO6bJiS+V6f3HZqB71hrZt6ymjF/kVDLEL03JC+nTIpayjRFuRbHv6mWS
A0vkl8CRV5OBy+mwLqxUyYfnuTm6PSFyA6qoaFfewKIJwPZFOpAEes5IHhCW850C
ZU5MvJ/dinWfaIV5KPcrgTMR0k7s2d1SQ1M8zCqfJBeMr4fRIapUTa/NjpU2w8HJ
y0B/cKtvrtEH12cFtoti0L1NDc/Bw6gajlGnXYUxuZwXSmgzG2JraFV9o4GOdnxx
xZuGJRUJe/TJrYqPTH1eTGHgWNLd/hGNt/ft2o5sZ/w/i+9DlkONvabuD1PktiZg
rDdgUvPD7RQXsEnb6/rtfZnVl41982HbTtEzeE+8a5m159UMKRCoE+r90VwU0Jp8
npgpJiATkwLaIxdW9Y+I2F1+OrJnH9RVvZ0OdCBwd0cDfo+MtLlxFKZoP8esnxfP
ZdRYGXqF9G+Uol6g5EKt13VooF0NzBG4u0L7WDVR2mCPNzR6m+e+XSiFLwI+fqr5
N6DO0AEjNeiZO8cLVnT6EEl7lUEl5lE+odjPjGHE5lWRitLxILXqggtiEsem7lwX
DKwDE5H6rWG3Lv8vkv07pR9CRqtS+foOxp/lkHIQbbNeQJC22pEupttXDzvZYUzm
wgk7SVSHSEYlVaL2O6FDnvzOw9TCemsMWyY/+GpG2yPxTIgyLyrObyozeAhSKzwf
GGhfHicMDgCkde+jTDDBaNQ6mTH3d09QviCN4+gsApbqYOlNDAwD7hsfPhWCmyF5
UQgtjMUSE1mm/dHFEONGXAo1SCK21AlgZ1pEh1ePtHT1SMBXbizqheM5sWmEWw5x
9YrOyTNBlRTOLaJa/ks+MIHr0Ydy/3M9KUX662DH6alNG2bOlaqYVx/g6xE6nSAH
WAiQOdJISJQDLFIG3BaBgeXzyYFruQj2izgd21Dq5pjwPJiCyVEtjqjNauPvnOFY
Tgce6arDJukltAnSYjmohq6PuKRYskGbriXo3AzJvNLrb2X8+GpFA9NcjquTO4/A
fMxSjLBNhvWTDnSGtPIln6jcK/e5SSXkej93UUjThyDi9BcRthMhroOSNEumsxw9
82IzJ1ZSQfnL3N99qmCRxVXmmEgJCtwE2JwOFNFHaxaIRFdUdPi8wm4lpsXp/0ZA
ZSrIUN0DAQ8UmC/uY/+5EJdE8Ls7bKwUi2J0AK8szBY8Jr3ItWtcONN6JVpPESx3
1JZTr8gk/pUrJeuQIwag7L4+YNUz2Vjq1H54QgKABl3R2xNomza7eUyNOrs/YLBM
L4NhUsrbYCcGYJLcI7HknSezq3q+biq6njJ19yez9Lwx6aA3rpEWHYJaQIs1siSc
68ueyfvQjkD3wdX6HcrQ5m8IaVFE+CQOQ8JsTrqg8vGH/A0wwU57Bj3Hft6wCGEO
xWIdOHQ3+P/4M6sVDpKupCDXL00darBu4i5a+p0XpwBtvZebhhuVGAHojvCXZBSf
qD+WtINx+Ep+C2Rzy80SFmN7mgw3el7y7VNfb1AV2eNoAE5W4OJQy26FD0PwLgvx
hr6ZCtUNaS+WxFbPIsCINo4MnTYS2Ddsf+WI5equsAyCxytyGwqsBcdTjC+649cP
LraAM0EdgWqZ+lrahOJDPbjIOuGS+87A2Vc+dLQhjjRuP1cDkSNkdEXGj8+HKiLS
CUqYftd3RodgXj3p+BAMWggsj1aHmgs2NS88T7UfKdIIBi5LV2gghd7jwqfYUDYC
2P7hjMkzwyK6BZ7Tx4HHKMjMQCdsRo2ikHtSFFIYgb5IWNNHuWH49m6kqOenTKA2
CNmrXUOU8r4ZGSfSXAOCHQV2JOKdkjo2INOExz9dqhgX4e0YQmF50ZPKDRyzEiD7
kcO87yrj90S+NelVrfsYVFZJyiCLL6IzEX3whEbVvLIiFL6nyG8tPE/YBXAlQxlg
UZ8jpq3r/jfewkxZeWq+m73UViqNmAcrRbQu0qrnvhIqWWL94LeBrrSz5ltCftOq
whBMCdpHaj4wvyb5msxmyn55CJm/7ms32bMdQfSgm7w7ndIK1bd3l2s8MuISvj1M
wLFrJ92XcHzUbsILmGbUy3K85cvurGhT2dm6DA0DnnwzX87f6Xs9YrFGJH4j/RmY
yTA0dl0oX8D2FbtrZFQ9eqH8NYoFbrwH5n5ZrNDGxQQROhKZkz+qGCgrvbqaqI/s
kYeQzTF1OP7xhci2Jp2tXw+Fnlxoi/eYE+8aROpwKXS1WcKmK4uMA/wI+saaen5e
jYuF1pRZOBz/IOKvm4h+IgOO/r4qTO4ovvIdFZu8p2tYs7jFXbJY1pQ3LvgwYEc7
kEjLdwQTMvGBhX46EQ33c9tHwkI6qGH4RBhj+ryjh17CoRcSMsNUvggDzpwrpoVV
9R/ieFZpAFiNYngMhCS8iHjRpOjzSqVQxuPrrAeKV6dolBB1Shsb512u8EXlC85D
U6UsRvOx+pvC1X4kg5inT9KrU4YMeYnNv6eXQYnHsMMZBYQL2py81bgIF62I9hll
XOuAcYdHfvMCR1ZRWG9dC/bAfkM5ps2j0NqiP1x6lo/a71rKgqrobbwSSdfuNLta
qGbAAp/1xgA2HgoeHefNNeZTVWmF3layzHZaQxE8O0sVwbpamNfkOiv37Ox4N7Pd
1wxuOIvqR6YRVPF3CUMoMyRIXa78SrFvIhRNkTwMfHYsrftAB4EIbHh5aK4Ky1bu
lCUJTYcTnXo7Rv5zaWZ5+vib97t4Xc5SPsqg2k6JYqvF1T/ceA4fe//wPRAD0NPV
lyw2QcuCSRdRvVOjJlCJqA+mRTkf+alNiddVj2LP8d8keao2SMTk7F+T4cp4cgJ/
2tq89wWPDErW5SpivZ8H7lQVLgfXh1a4GMjyY3OK/kMG+N9PzfQyGNtqS2RKkgnq
Y+J8oqICYZf4Vx4n8+BiUFU0Ks7ZtZeJJynUSVgkpb74XN4tdtFJRhaxlSnaRgJl
RojiBsOWUfG2XA8VjExl5RQe9jHDSZHbCsNMvOJHYYTmxwfmFfCdLLrZyBt4kF6h
A99wlEzD/ybdSr1DUf+bsGbLfARv4qNogGGtG+Z6zm04qDbgqGCkp5x9oMhnwp6x
KFVIVys46Ckl0p2mFZUPBky8eMJUNeRNZPrj6x2JqE3JspjAJvJtJH7PNsn2rsDO
EdE8BgLb6fGj2HncgpOgt0jV5+DCE1TGmrHXc3i3FC+kKVZuWpHenZMVAxTcXQkE
CH2UKSrF07kGVZdspricIgYuQku52ccX5V6cCFy60hR/jQdIq/Bwk+6HJLwcibE3
GwJetYT/emOKWCe7aVs0Dx7BHdF9FkftLNR2e3lZqNaHuGwe4Y2XpQbnVe7YW5MK
nmeSpmKysGzITcjPBlf4kSv25q/TKZJmUTVyTJ7b/3T1qEoFFBzonlX4ND1TNJAg
7LVHWPNTdUtiqBkF+bEtT/lG+Ts94IotfKa6CdmY6Xz/dvwQdiDRlhj+wOYxBtVP
VBaklsHzxJG78qcoC1AxngicAkqMq1HQsXcmx+XVUocdTHJZggBwESrp29U7E4g3
rHff3C3Ae84kg2skNqR0k3T50rqZaZGjniLPHuRI1vg8zRsFW6UOZd9ex3CNVdvd
D0oZR2U2HIxqzJjmGEFtd+Z8q71qH8WntooC1qVe92lmgiL0DT0XxvJmZ0RTQXlS
c0mmP3yeIaaN2BtbWZiRdvEKzbgDCanZPcMWTrmyx7Xr0CxIXwIG5icvIOAC7uhu
BbTuree5xmVap/pgaeIXfxqmdVZBHtlTiorccTy9vBRhbajrszBWNmzOIDNQxVCB
vfiLtha+5e29nmjU9XH+UP/ujbMjHjy3s3QburTxLegqQCu5bYvmd3R9MM9uZ1vT
HPRx6EcCosVeL8NQ2d/kU5/0i7a3ukJ8Bro82hmIBHvjtfW3Vtl0CRNiwNrJDYo3
Jmdc4Yf7JQdlfEnNoKgL78+QMnea1pcClojS6ExsM0t9NQff82G/6PN9A44fUeAT
sAuSFwNRGZ4P8wufpK0ehA7dRuk3WZCyq5j3BMBnY6d84tQbLzX/VBmgaCxpxrck
orJ5/5cYkGlMzxt4je1Fdi5OkM/ZuOGVf/+JOl92XUHEA3UMWmkabMUKg2oZbk5g
knFy9fozjQyr3zXCaJz9cFrmi12IHskOI1mI0uUzrpPhxQKL6LFI2e566ieP2ga1
rOAc97wIOUWnjY+Rp5BUToilYNqb0pVTjWOaalU5Gn5znpRVv8Wvf4HzsY4Ai2DU
0zewpI7Kde1NeKdWytH6WNS+Nwe0+YBxrM6KsQS3K8UhexXsroe6BnftXfDRbkPi
7I5LsjMkQCusjHm1QAAmQ0ciNm4sXFPdvfZgYXY/f0QqMu3Yd9Vk7q80FyQe5ikK
JyudZTAfLH8joMj42dmgi4JOmMbzA47vs/3MdiLWSiz3LFnMnvpfqBExZPr7rmYf
rydafnHJRYdjkq5tCgB+K9BneEE585ZViKw99N5cPGEwAF1kbCKqmQoAf0g0gGtc
yaaaGIvIf5UwGMCEpuQXnANHqHIV/JwF6fZyQoxESYgsJ67CMPOPXUk44grZkGTe
EjN8iebyCSZjblYMJ7jXgYlH6JAUC2PuluS+CNrEoKXm/NKTzKbG0qBESLZ3ovvi
R3nDoG7AKhLMRFI461uVcr2OUtdsf9iXZZYow5J158vbJBuRlvdrICK8SGrml7Ds
pME4Kwu5SUWED8h+MNSAhnhkOnhdIjEo7pxGVDREQbO68bPL6S2i9Dkz6fQiz/xC
wUFGAWmVrrD6exmp1CtpD5ZM6uGRvfLs+Q7bjE1UYpc8ZhQ2BiHA3NY2DXSAKVsl
ExP2BL9xkKhACg++4nEk4y9KQnkZEyuZr9vY7dMplzIuL7pFoGD7coMprS8gmE9o
+LbaEHJ5qAxnzpj0sAz+BrCVbiW0BVC4Dwh1IDDdY3uSw7bVRqtkH/v61VuXZzyO
ys6ezwcAotB15GXdo9N+8sfE4z0+UBVVVSHY76Ki9+XXdmL4SIuE8HXFgrt9elPP
TxAoFkAa+nokERegd7kIQAy4SGBPRXQjKNOq4kEJXpTucPCCt6OJw3M8xbYginlc
7Ut/lIPIfKD/qyuPPT5c67pjTQ9mbGO96ZcVU7rxYnzRSGnMiKMFUsiocyX5yuen
qzeqC3qyqrBLdFWGOiiQAgCyts7F+fZfmQCwo16VB3Hpnr61IfebTXkI3jw6orX4
BMo5PLBhFHj/s1wbYFnlaTRBAMGDhx5AI2HXJ4v0mvVOaSYT7+BYzR1nW1DGtsTW
nmqAsja1rQPXc6Yw3BfKcs8no3r5c+j+M4MmJjNkncVvc6be02tF7oJlI1U865Ab
wlksBfr25r63QGbAT+VD914HqgOpuy9bThIeDzleZCBD2HH/k3edJlxqxb20u0At
fiqLXa1CliMjvx5XG/ZB3RFnTnz6LMY15RqV/DysYhl9QQl8HBVckk/9V1PUTj0e
Whkh7yA3LdNRKK4/lpEBTpETqEBxEmYEvKqZ/dCUNTsFo9Jv6mhYh/s239T5LY7v
YAry5ZZ1/UcAPYk+u3tBDoJih8UDEvaylRITs2u0w4mfwCs/gFneSzZIWU6Xe+NO
jhXkA3u9WrA+i0JE61v0WPsTU4r6lg6h4iQt+1mGW2dcK5W2zqgLB2GlE8pDQrlP
y9Jbm+E13JHIyYeQQnuLnrr623EwoKOKoO5ZH+uqL0J4xzvelbrtZuq/uZAjej8u
MCPvG8h0tRXKA5gnDL+oYeATUWkteKqTpVxec33K+D3lq+swL5EGfAGl59BwON+Q
NlbVFUb/ZvOYDImLj3yYzOqQ3cNeiG4KES2pQvRDxSrwIL0DLdIly4xmNffyKffB
nM45gV4DD0Pby/ADKITUQlhwlY8T9FSsl1NqPYAdIgTIEr+JuJaMNGPMbL/AJb2F
Vr6V9QsaD4vMnjlwNlAoZK1O4z4VJOVfF0omI0cKoZDlgz+IpceAisWxQAYNldtL
8uSjE/Pywjpzbv97/eYftdAbmb6ZiAzwt+xV3A56wwTqHZLeCArS0c2AAyOibFxv
kcsZpcErA9fPlrg4tBEjTcQrCNEYEojpbcxPd1eoyEOkBnJ6MHHX8oydsuJKqB/+
QwaNVrkFxV8G2fjS6qdBDZDSM4ms+axq6ZJnmvH0RJdEWpXaj1UwfpGSAWwptqQG
twxYgVmdaIt0F59xeU4SmgwttR1dt7I6oR963TcvGpt5v87myTjdGokX3DaEZIzu
X7FiIHktIbrCrg4Ap6WzteeC6Zx79jQ7JbrEWjnwh5XTWtj0trw899d8yIBA6AGh
SY1g/5rIKzelzGN1uTddI10jg2NwNCoZbySaeeGuLT3xXMEyYsjE02piPhQz8U8g
nZNlopD7k6PerMvFiO+/IHjH5TIdDzy/UuGyDpw239re3YBovPQPixhomYyWZaHL
RdRTU0OlSVmaPeggadyYZ/Wg1Yh7pzIdY/an2jkOHK6LsOMQ/2I2kEjOi9BtC6m/
Fcn5TKrKDQuwyN+MZ7qrBQascKuXL3GUh4fcnIBanHU2hob9tOUGOsZl0yMaqff/
VGiy3Pt14Rdm0QNVqeRDtzIU2XnZ3yPVqFz6RQmB0T+YsI9mc6e15bdJMIdAyTgi
e6OW2Biafe5wA1kCJTIOE4ILsunwovTSmO0c7on8BYgB7eC2zkxd7APLTfIK8Q9u
LoHTDvgFxNDqlECEVf8sNSc8vC3jwAjPaKq0jHNWlOmIGC4BlcS88yTk7XsDOfVB
Gy+1fiouR7L1bGln8LThdUc4zstGl34FhLLnUVWe8KHA7OiE/PuWd2sGO8Gms01W
8bPF4kKZaoxFkRFikmAev+Sp9BIbPeYjTpLM13UXGAKFzOohEJz0Dwo+Uze6CNzB
E4M0FIxiU5hQ1txaJhXSXekIl17RMNyhi6zFi9lIdZYj+fAy0pmTvuVLRwzZEMcP
E8NJkflsUUOB+pGwlLXmAxCEYWk/O3eV5YhEgQ2drUHsAPTy2YTMZg4rCR2omF/K
+QpvrJW2bsVjnDdjpvMAhLKQYrP38qJrqgEuPsHv/RKK13opgkGHv5ep2Wx+lVsx
kTG1G67b6tLVj9R6u8xpeiHLYGeojUDkuE7V/vtS/VnUSlTBaKTTT1GkZky/+sxU
VmUQArbhknTgdQ2ax95zT7sQkWv/JmpAvC4IGXH8/W3HVLy5QavMal2e6mBLjn43
nwV00WgR6WOqVWPqsXrVbpDOw4nVU8i2ZA+FkQitRd+rnlmCZES6TyU9cgB8HG9r
nEfrpoga0s7GW8+SpPzGMFzZ7z+3wJdvGPul2lOeO3Dr5UWUs9C6JB66qzJB3SFc
YFWtdxFC/tJ8ujnvy0TJG9dfm0rkYznqej4IMJvI/rjqgn07ZHDCI1tMsvq7LOpY
Mu9/ve7oRiNhQ5r6xei+J0hkgML4M21wpu8Wt4nfD8bddfIZaqIsQxbZHdqswlKv
yvG1ruyGyqyJdZ/UoOWrudlS4vYjXgHWuFojVeurnhSj4EWk4yEYk0Nvo35UdloV
wuXqXPzMq4DDvPZnjA9S2q0oCqIyifdWcqqJAhrs7YfTgkLzaVT3MRT18LfSTTQx
WdBmc/Ih08kpVfzk56SUjHSXVahJatns9+PIvObmihWV0ALSNzcP319KJV+Ahvxg
99vAvP0kqBlwizpICc4RvAdumhD6RfnBhpX3WoPCqbgrsjIVvNUectsvMnDEG/sy
Eb+5R+GX/8lJ29ckimYrRtwS/hlEv+whSm7lbweNGPBm1XwkNhtFSQGN6hgA64nb
/5XX1XHtiDwZ9lv9mRoFxR+JLa527UwVnau8PRGFtlL+kcCiyZG3mkZl9Ui4FjaD
ABCwfYRyRaNwhQlH+qcAjHDnL96MaPBPalXPedMSLrT+kuXNBcqY6ezPY1IPpwfW
Xfd+37xGr2GsRlezUp0xtnHvEz0rODj9qtVd4lb5ggnuBWBbSX/gO9RNOHT7/IPA
fzuvgYSKnqQLA6ag5wkIlqhWbRzHlBa/2/h/QczD9rk3UE7yTM+4H/6INvyMD2KH
ALd03NCwzPJ5Hde8A5VrHP0VeiWEW4fG9WRqAJwexEe1lgQjH+eIBRx0Cs3T7LUl
+38qbDMc8sopweH33rEfiSIlqAo2orlz3CY0NXqXXBNGlD/mf+IOqiCiveBNINyI
efmLhHa0gscDNBde+ZscLVghtc6n9xBXDs1a2+PrJBXatvlhgAgbvJO2HcEqFLzE
msqHR7fEWdTBp0hKYOYIIOuiRNVCi2tu7+KcVW69AFksIA2pofRFVtnrhWubpMYz
cQe//XWqXBcktnCcoXCF2iFI0TQv+s1DkZB53HKabF6dNMJC3lwQThSWpUVAt4/f
kyATrStP5YGxAPBYspQ/1MuVwn5ps8n4C+bdbrU4FTHlNpaORZY4wEszJ8lvSLeM
d7g/q1x3nX7sNEfGtyFx/SuwsBhhogZLcW6RCXuzg5rbef5Sek72bj/Mk2s6ATlG
88yTugrKKjf12op5suALmRDq5SkMDWy6T1Czq2pyTXgVxLfotIlZsTI5cEUHAcbW
Vl8lknnggRyPDRaCWe/96roROPXmxQBPt9wsULPIGg9pmidhFy6MoGVuVFVisnuj
gFwckxNipyT/wc1pHqsBTNyPlenrJnDaH28P3+MzewRIKWw1ARAtwT84E7D56ghf
FXcssEvKkj5x5FnWRNxghqyORxxyKAxPEOR2N1yxvrr3yB+sbgDrFtmxEAU4UZEn
pv9Jl9NdDC60VScLoBl/rtFas33nNj6m0835UyZe0GufvMKteZbKC84cnnSdjjcl
zHvBY1SqhqsgKsArkVU+fZFbcyArBDG7C1gKIz6A5pUx/XDX2PGWoqjNIlfYWfyk
fCtCR3K3HLQjf8BN56ZemhvVeCYmqmYtcXZqA7G9KJ9/4MzSrrAFbSMJNqYP/ULZ
twNdBuXLxGno4/IXFjbS58e6LUNfeV0VVCGjCf16mTQj2Z2H76nNAdRHWxftI7Aq
fRBZj/2QSaEXaBr9TlL1doVxw9vF64z75oyONVAUK8fmqu4lCZXENQVqs5F9AXhp
cfkd66HAPufPzUggyY2KtA+eNVWa/C+CqQaSaSc91R6frg20FmF5g42T4n3b0/KH
nR2wbMrYjkH2IwPvRoi1gJqRX8b7OrEmfHRx447zUSY8contxPpdP38mzdf6PIxV
TyuZHF4lAhF3KtC9zX4ZER70nQE717c+R+crdpw4tlzkGbVOukbTcl/8+/iaDBNT
MFbgSis9NBt0/opi18s+yreDoBqeYnqg7rFpDUPF6VWQXfkEJeG0Zb7LB3w9F1R3
+GYpV3ItadRmnEYM4xOYdkWlV0yz5ZaVFVgBZFFMtVSdvPmfTTiLI9J0N1Ogs/al
QQh0tPV6uoaDp6a0I4Ark2Ty/COOQbHDABvZNjV3JLwSMF4T414I+Lkp7aVN/3Oo
1EVA32hHTgvnizoxbX1z7C+kbB6TPpScM8fZVFRKe8eM4f3kV7tKt0G/u6/sntaz
YskkPI9vftLRVpPU/fQUtdXJ2t6LmAXAJnBv83SKft1W0LvdeaWVG4QcSUCXZwCa
I+aQ6OZTlwxpWw8Xd3EUbEY/Pu0QYNHdZ5zUT2gaes9LmwxxnCWTVHqRs/hphkL+
RiLG39jwjPn9aSRHGW/BMyYqyN6fNy/pnqPO4kk8F/7A/fk1jtKtjzu5Br/JJrU6
NiU07tJrIs+yVsa8P1JqLbHeXMTe3c7VzkJvG4exq4TsC3NOlsumw7uYMezuCu6j
opaAV2Yi1ZpsHav38XHPJs6FbsL/IuFzr2Fsc3jd2oK0kFFygIvgP4hWiggIJWmK
6uPZXE3eHZBURAWDyk9gNUFXrNdpvqv/a0oC97nzJhri9kDg0vI6WXbEPh126ukQ
kOHSVsjAY/kLccup8qa766CyewsqHUopGiSN9tOEm0/1VbWoBfQHL/k2I64HRQ5k
qCqNopq11PIOLzva+f83MpysCmkWQZmQyhpGgjfQ7Dzzz83SIe4e5tk0PeO+phGS
2nQ1YYMX3BfJ960ZEC2qWET9aqNqGSSIT2xa2OCEVtjyUEaSaUMsgj+hFo/gPLfH
5DlsGE6Dtvpe0pdciQw8+F7VEAz2Bdc2dvb0GdFlSaABX/rnwSliqb02OMffnkGv
wtbZjNNZgCMQ+9kJbW34jZ/vS2bxUOOE895N9S69btEQ2DZy/ZY9nJJ/yD5kHx1G
CRW31Js2n1VdrRVTbizjxFWEeMjnyp0B+8mlbDNkJnxkyjEsts5D9k9cFX/RM/mJ
CHscdE9yy3w+ayE5BI6qiC06ZV3Me3R1/PjzmLWfLT4XlGH4XENnqbYhcFsstmQC
T34dkenjObiBgFq5DLnkLr4YLwicbKxaikgdQdsgZrelYnFUntkv30dvr991NnHd
wqhn+/eUWJKd+AfUN77hGHJVHMX7xuKWpE1BokZVmpR8kb6nKatQFNuJjBcZbqLD
Sej3yaIkPMHmJLdH144rQ+wjAUQ901Nk39OOfziY4YWf53RbHdFPoPhQG4wCZecp
gyf+mxUStce9VhBYlMmnfrGg2Kj8jWZRn0h/CHJviiZahc4FPTupDHiaPwh37hSF
ylnnUe20RcP9n8SrPwtaoF5LPTTK/8wdmyPVFF/7g4DFwK/jhs38kT1trsRAzJaM
FQ7DsUygYB5iEdw9B4VrB0W8ml8tdH5phgtkcprIRjSFK0wRuOtdKKhNZLlm6gMm
V83hSqNQ6NoEjhEluZeDLAA7moVotzqHj76OWqVcyYrCF7x9Jd97vV4e89nk8BAV
6ivmBwbohMDBcngqH0PdzeoHTv+JvYH45N+k/EB2NIU5/u5ur44lZua0G8wmIzq7
luFqQa940j2yVt+S61KcqmP/Bs8v+TKdZpWuHdWZ+vCfYJWdm3odNoqw3wH0Ably
lggC314k/O/D+oNlX+xnxzqxLiBm9zkFUw4/onQnErkNvTOVgbQdSRJIFQsGBW9z
3PNgIzFhkpPxxxa1k3Moxy++tAvtohll1RUpXXIPi+HkRz3GRM9F7twoWTspLd/O
/ei23ISraNnO68aJXNuB/OSBulpeFlvul2Lp6iGiTL+H+Ze6GRsEjL615I+81TC2
9NXuYNSyNxlLBa9YymNPQMWvxht/IQWB5UvX7z+XAQe2W3Fzp/JgDaTM3/h8+4zm
bTws0FejmG/xvkl6eVpy91H3ODDfF6ZH2G4Fx67CwnN6Pr+JPep/yfs08lwEDsiu
xS0RCFmEWC7NmIZta4wG46QURQ8YjsBjhCYdjd/gRJOiLQSv33922lW3D8mcctbd
75V3AFd3/eT1/1Y0f4CF69gwSActSOfjpGU8N2EBoZumy/e2m6WFtRnCnAuG6ATy
1jSmfSGDB1FX3BtKbgRDFp5y8lx7izxiATJYJ+949dKVF0NygkznF47I3Wg5MPn+
RnwUgTjzsq5uMEe38XULze5vJ6ts1lTKFZpNfFyA5tURVeOHMM5ixfuDIGxvWiOa
3kF9ma/MWWzQbLDTAXwYUzzHzHcdIveDqkWBYC+H8kaFs2JmGhiDXg8Kdov+AQq6
RV2u5Ajco1tJRLvu8/RFMtjZr7nER218fmQf/hKhzzHbyAoQTDQLJHhbYS16eoCU
/vf68zddGl0UevAcSxCJSnSt7b5kFlWX5wfP1X6evi/E1U7YvWcXm7IFFdwFAqf6
2RyZhIOhhsYo9kKzY2a743dNU7qQQ1B0yb5/blJx9IlodEhnUDJ8qFG3LuXYcwJv
sPYt8C9gtCw94GKTyHTHqRqznSX3F60n7lP0+kAE5+o1FEyjVBqWqxnP5ElH2oF/
IELLVWsMBd/UXkQ7HidsZTqw4cZamTb+yHR0oVsfAMW7Xu/9SCY/9rUFUFVB1k0Y
BkZlHOuU3v5f5fJlV55YYol3WImjq5sQF7n8CK4koziSZz10hXBzbOQUpd1kHXLy
GStEl3CLA8pHmXbczBlGgqeOouZufEwi39BA9Gir07ESQzcVtMKNwZH60zxWOroS
Sdv7uTgCn59/TmLBRNnVV90CQ4TsFL0tvqV/L04+ZbruFxXOh1tQiLDqksN/POsl
G0Ug3OEzfIy6eXJDPy6zNdx0FTO2qwNo1b0JxkjKSGsOAfs2OTulAaU1DfgGSy6I
xjz6Win9D39hAMsgDFyyIWMqU8XpsEtYV9cW9DWAtNZaCRCix3RKkdaiqJbbQmRl
tWllCQ3Auq+uENsK/XmjMLlWPcW1zpuiAuy3RSMKvtd9MfB+3EZnwJgiQoev5Qdz
EfvjYOCmwXDUK3f5TtVxmR5q9I38zTRDnqfeYCfw/6O+9nCEx696Ym6H1e+zDMfb
o3TKgPKYeuN1UsdhfvZtBlT9hmNAMyszbKuNb5kd98GZxBrICf9arXTRL8SwM5vR
P7ACmATlYf5ODpr3Fp7E+e+a5Pycw02aYJd75Ip3WPqWBMlnNq08GyOBJStRjIos
ohtKwqjkK7RrgsVj4S8dR/Jeyg3gdEqdE4oXl193x69r+v7sjEKhEmrQyX+KZ9eb
IO9q4fq6RxclCLWvCZPQenUTfCmzaZLJUhaITK03DaJFbESCuvi2oY/otQEEcPPg
sJZQ4soXDpUoo8YdxyTRPBDgygPFLDjo0NLHjtqHIUVww/4T+EYd5s9VGqGKzHt5
KBoYfz9a5ycLDrzcPDwW8JdgxIzjuMF1hj8xobLQpsbi4djMxGXx4KNzE49JNwWG
4JxM3fKmc1jjIT1aCVfIPJi3CbW+A7fAWYPezJIfpiKZNEOumHkTRlQHYfxVTLXw
ljINUqEG15j3jv8faEhdZo/CLOPysDxouA3KSVnTQ4RpCn+PqzrY/NFUUcRHF1js
g9orGfqTmfhOlZXxIbjqUIwoRYo9aaHS5VbaYmGZ2ddpoYak0cHYsJFRQEwyfJVP
mKqmkhOyen7T75ua59heaV8TT3tifM4FCYyo+jCdlK1846Vqnc0Z9CbNyN7rGUAQ
DKac1ZO2HxjerczJCH5ooCU7iUOZ3rBjz87JGB5X96DQHnN2Y7gdmVo2HEqYEvEI
i/14AzAkm/b/yvxOEK46WGU1UILCJ8dSxf6KNv4ID3z4a33L6oP9no3+35IPqxL1
PZNrxXBCvlQYuXNq+QNnXbK0eoZAcO+xd8PXJkbjM4J+eUryam43MuqHqI9GMDTx
RMejmlV/5pIFK3v9DDOiz2uB1Ps3tBbjjzHh02FRtvvWJbhsb1/lY1eLBdt+RIAH
n841wTIC2mUaiCVdACCmRoQQNT2rA1ndOL9hovNXpfq/+Pd7vT2i1ggFS0Vym1yo
N53J4mDb5l+uVZwWCJTQiDgzfVcR78rS25Bgk0bCYIF/wrs5Virb94M41tjljSga
4DM1Y1tTlLallsOrlRLaTSd7eq/uxDzPEjR7dLmlzNziCGjTjMgmH9qnB0AKVvBJ
WR5GPDRv8WC7+4DvYRFNYhpDN7h2MAWIA3czxUZJ49CMAAqK3qaR9TwsJwEoGqab
BPLMhkiohojzbHwrgdbSnlfqEbd5yHsXd8aoId2K4M/5bDNjulEgKUI4cHDPlo9x
XuAUchvIwoRT+RrikkcdnSVeEwFWWwfxea6q1RdXSxxqDABa7wfNL//PNOObzA0H
glLS6EheTJgPiocxEJdw+oaz3u7Vshul39mswEw0Ci+nXigVAxCZ6IQL+pVRdWTl
+CRg0IE/bgmZLCpqPxqrRLG6+8zZ3hYPa47ptl5GO0oFuo1bEi5DOu5bzbWsBS+g
yAAqO21HsLm4aoV1HGFxoXhqwvAfHhijtLIEWS5+PkpGpWEDXxPrriE7OymG8EO3
vEiVk5bxzMn67ZNUTxc8/LIP1UFx+2P1HGtnZEasrThEq7REQwJ6KJeh4h3PiglT
+db8RI7y73zmfSyT7Q011cv/SJ84rAeK0P26GN3bPfhMJ+JgHPzI09eIBQFOmXcO
lZ7knGzS8Nr/v6HbRooNLVYhQJ/Yk2mjUAP3woVRIj7H61Pw65x2QxRVPNEIzU/Z
BhYhGStUbcFBlLkKiMTdxtK9OVOOVjGMeWD/4+jPCOJzgYhZ9dC3fQEpy23UzoBV
5+hQqdGfNZ99SSKV+fQSTFJbIcmdWE3XyBUXx4dmRHBbMHkpw7O4rHqN3nruzl5a
Yig1TvoD6lOgprSg0j8uyQiJfvlf6Celc6YOLAC8DMvC1aOdjMnRDUMVS8eRJXqE
sXY4Vk/HMPBGoeWbWiwdrKiLlKgW73pFL6ZcUNof85sPAiHxvMfGrHW3zPV0b6rg
Z+zOd0a9q1/raTjJtZGrNnM5fTb5uvYPeCBXF2shpAfNER1e5wr3cfxmzFdVPOia
e2wfQZevBha/TgmMl/mSw9Rt3DQcc2OFBIZJPpBjQ1kapq4aNQmME4paBEUE3c5g
t9XbLhN9GcE/W9J3b3mGjSp0n4WQkuGpdRV7kEgV2R6z3e9SnvBXnWcBDyjkOzXi
j6RMkCXq2hSeohzA9GCjX80Q9P7Zb7SGf5AVqWoCOEEG4CK19jE3mhAEZM8rB2/b
/xg51A8lfrVWN+69STgYJTXt/cgrz/wHGosqLEEtxdHuVhbs1KF39sqCzO2KBbQw
WmwVxGkO+74jH+UdGa/HXmFgxvU+7VSr9jj5R/RtwFF8/HNpLaZkoM5+kWFBnuX1
2I5Ko0xB4H67e9Z76mKszrN4VviK3eIemLHKeIJOoKUa3o6l1L9qhK941S9NrU6G
Ulp3eaOS45l7DQL7tXaBvAjVT9VrJAyOyMA+dUTJkdWtXpZfLGgv5ChSwUC8H0De
FJqjsmGR5iNng/GMBkuaJxpmhFPO4ysAxqT/hLeL1tPYIp4IjJbEYmmdPc2kW9Cy
Z2HhYBbo7Ar8Gxk17dcTblc7WT0pXMDp8wQpuq4V5leW2frGp2GuNtu1mxSByJHM
w2Vu3G1cZ4fvptgT9LtjX5JardSHvoehME9MuNJLqnGCmtLPVmzealZxpGejdYpf
zuGVc5KgeFBSHH3bRyJMPOu+WO/nAKtboc8196q9XfXeqDqXRsoIG0dEFhG7EDLz
eZ18xD3TusyO1028d9kFGGAz0UPXSa5hgcaiMCJdqhMMEB3SLu9xGH5M6w9cIQaz
VgHcLrM/kas6yhvLgZ6L0jXPpW9PCq+pZIlkjqJGrgbpERea01WdrYWKoCVhIUnN
6CZn7YTBSUubqDwxscikdlmYi2x1fRJ+zF0hcKHTGd6Z6Se4OetDdzar8qBRZXJt
z3iF7tdFOP9bAlGBixmOBIlt/xLttAchhOZJzx0GKc++OEZjIxk5YbBTdB5LRzPc
RbxLAg4lxF9Opb9DDwcjl6vIE5JY0ioCEXP0N19fF4LLZLx5RBr5cW5W/3vgnRQc
MArjvb58SmFoG+FSjiTmoNgsoKszxECdGYDqBvvvYM9y8FWqw6EiJpxLYSiXgv1I
UDUFpXqkxmnYY5JQlZi8T2OzQXgzkfwmuYiiEZ5UtPAi/YFbHg12GpFE/CCSauzq
Ymnh1BTYmhJBk6vznSo/Bw68cdo62XtIvL0yUON7Q8xI0ttLhT9LM8NXRqY6Dr6N
S5cDvE7GFfvra2uO7TnaRCzrn+v2Z6EkCJT4Y1WO1HUpIkiNF5/KJtS2DJwNQRx1
pFf4ZFRT8LCFmC/jQUCozR7mxBbslJr5uZRAf+vMEDEWIqJK7v7MVcK0rSQcJ8Px
kfYC9U2kMNnWhhtYNIVff4VE66GEQehy8IigHYPyocmKWVhVMPxCxZQgCb/KlJ8o
iwbVNIgxfSn/kMK25LmBuprSRYoBxKTi35rttBi/xVVOHjqWclGSpfJhdKCllx/+
dyFYsJaRX6mjQ5fyLFhK9IvWE0d8D55hWr+FuI3X+Kqnd9gHKd4XBD8fWJSo5u3S
MB/6Ix7XwvcGL9Si7XWgO+TY7FalvEHP50VtHOQBWKg2XS+N3e/BVtBmiERlUSrQ
XOg1QV/hm+w0kSpUZi95DSlQBZV4F84npl40hpIZg+++WBR9sa041TC1tFdvXKvz
iLyhmZJl2Bwm/W8/7HfDRhlBo4ynQD+lM/Gke1+i/ttaqzqHXlMo2E3r5hvej6Vl
3yL4+wDSi/Ji1xgnixo+ZN9vrtFIbUn/TwgzxvimxxoZIAYWR6iPon6RKJVjHS5O
txP2YjrdyjH57W0rpiBwT2Cd4Tn3TM2+fLY2QIj2ZCFUyrkTAedX7Ob8NtV91Zp4
/YkWCqnXbh96TrPzH4CL2b6jpXhk0EnQhyfZkGpvqvAn7tepLPch8Sa0mCPip1D8
4ntc91yrMVYNCS7BDKRHBYDq5Lptc7JLDIKZcysxQI3NRGawfC4YkL40HbeaHntE
ZpVsIO4JpEce6P5dehi+sHVMXCwCTJJ6D7QEZamrDS8R64WvS6kKcm2B0efTOxzk
UGxNn2PqSIlMm3Ivids2szqDTsXpJKq/aVNJ0cwq7oXTOXrB8V0jefBL/ez7g4Si
+TQr2sRAmJasXcFotjqTtWW41Frpiphadk+ii+P4UoeA8UnvxcOsFW8Lh2p0/jSJ
kI51bEC1nivU5o6XYEBxfdc2XnoTqvLFFdOoITK0BcpBr7Nj4JmZq2GRgzc6ddBz
bdzT44j9I15R5VGb/GVbkhQAnzJnz2CueRnQjfDx6gxbww4rLf2X507KbkJZyzHa
QuPLdCiYIih8VCRsdvU5N9WbV73EFPs0zG+j8EpPiK7RAGjLCQOtwHGaGHkQSOhT
WzFXPw5eG6shw1Sb6eMDWcN5Bf13xPKSMfskt+Eh0FBtgsnDV06z+8VKnxtNuPLM
nuQkybuiiBdkPLmbdUEtTrzbP5OBuDuZQ2VHp2pU5CsgeMMqHArW+efKIRfbRtE3
DQbIjOUUUmvH6DvAfZEBxnmoZ/CjYRD5av/NuO0Tv9Lxts7cjXP1PUMPGISHPcX9
S2hPG/ueykzS4EaSfTRGJW3G+hPp+shLKPPvT1bGJDS+11JWXqO0XXb8C624dUrA
Jai/k777TPOMlRpx3Zmo6e0rTg3Tz756QTgnhAUY6vCGhyijrKJK4Tr4T2LUQzKt
2tz23/VCc0f2mrE1tG/N5wJ+Xlj8V8EaDnHDI+ximnAFdmvgTV5gzRfOQUMSJI3G
7FqM2wKiaxb+nFblFMCJzJlzeuFD8BXpNKiMJimSZJuMybGrnqGbZBgnzCvZbz8W
8CMRrdcqGTl82VLek7NN3uMIWWbspV+XAIPcCTuWS5p6gRLvncq1LF2Rhd3J2hqT
9pjIsrT5imZQ39nuyj1W7DeIqeoVq3yKEGONCq0J/0uOM2HSZIbgRQmtLxrtwhEb
Jtr4KRuuenklEyYIRIr0pK7ioDMDxRb80tiLqvU+BtZuyQ/vC5maDiOHtP1iP1HR
v5wcK1I/GYghEN0I6ArZ8EY4rb0Dt8F7ru2qkdrUeas9vqGvodtkiq5ehWen2mdi
wnvyE672tef4PPQ0JDJha3cYIJ11LwGi7zZ7WaAjzmWox0y4A5HOlURIXr+6J1/x
2p0ZKSW0ySsdjTIhiU0At+FSrPvftLYP76iQ9FYiD58j8f4XG70OanqAhesFHGgo
oUpO1oRMygI1J5UIZq7Eh2oeu4JVw1pw/D10Srv3f/0NEmIAM3gydmtkdFwiIEQ/
KcR7U20V2AlO6P4211ulk3ivelTrZlM2J0XEUVlbgZhgLQYe/Q8/1Q51qHyAtmvz
aA4vbp8xH8+/S7yhFLLDbbHwhxyAq1c1XPI2WZWhlimkeYPRgLXbNrfaVYqWC/kg
Jjrkbg18G27ne+8MMagIQHk/JSk4E54/o8207jVcVwmSPt+JNLm/tkJJ5Jt/FYli
XTvIQbu/XrWvzID/OkLSDivhZLdANcpG9/9nlvqh19p/rLGeSwo6dobUjavN/Xcy
G3AvqXNKHcTtUqr5jrUtmMaTlgFPvujiB6ffEYoddAwcH9VPaedUKfdIBWBTjcIT
A1AK+z/DgExqU64HdwHyXxzsLa+hSL56dnnuLkDvZqJQWCrhnZWtj7itFwLkAdfM
Jwcuq0G+n3XEYN41Wa3nN24+eEGAe9GU/z7pBb8ESuAB3B/XsDemcwCdRRixKkGy
o4GtNMJC2sR7IdQl/qEwo+CrJBSeLNIiTLLe6wSlgVZDJX6kaKognTuTjEMDlilI
NYYURPIBmh7EHcYTFsCf3GdJBWJpyu3tFeCw2HOjR8VgeXzLfrj5qyvbgemXwxfl
eet0WZ5m6IjwzbP8khE6LUMMR+bpEeSF9rj7FKG0si6yK7CH6tUfYS8Es/v8mANv
oBG8gH2r3S5Kao6DciTXU5GEPuQwcjCoKgP6ElfeMNF3rCX3mjw1pGq6Et8h7jAA
mw/CXlYs2InQ+SOe8ny1TUToVCdkq9WP3x0ZUIfRXeat9u6DWsdGF5vhzVxy6Qe/
SRY0321Xms8Y9YPaqKLHtQ5TolVms91B9VcvoQoedbJLsiHEI9AyegKDZ2HX937i
EjA9CHpmh64pGCJi0/19xiC1Av6oPc7pMpgkldOvYtc2cGnhdPgSiZjdtKLBC6Uz
V78mJTucCnS6oQOg7wzMaPvitiPUf3bpgeCNnvJ88WTURGuJIO68SGN+Iku5swO2
Kgy52UlwVhvwsSuGEFXVakokQjaGrtPlmg8yiGCq6EwELUp5dHYiuJ9WSB3A+cr3
ZHDmC7bSqVtbXGJNWXjyJNgV12Ag4ANtePj9GHgDerrqOC5RZioF9Hb3a11fmQLD
g3cGBHt6zT+nDlTol3vzE0U/9YH0HA62Fx+t3a8ki0PZ/9SeOihCIs6l9RZnQ6OI
aBHjtUI4hGMAa9LEhh4rApHGTn1RI5ovHqNTD2ghXgb4tWX7Y2JqQoinNCiMInbo
5/d2zpoBT+USyRrJoSj9ofJy4fJww8o89etkapg1gEaT063nRk7Uh8AbLnK0IPOr
fvWbzr+lFF3zNd52nhbDp3K3+e7TTiNM4F8yPuLR75hQrDMoUw4HP9gX+LWygH0v
MdtcPsKzJqRnCzXV1S/wr/PO6rXUG2LiVreCwGW4yUkLlBZcJQ3cneJ+J7t/OsmS
BO1layUxbaPIJvEHXXcq08/Yvi5bFVMUmqEkkiIa1r253dsh6TkQFsUzopRfVvYP
RSExOac9nON6kQGBGg1tZsS9vpIuMvDpAOXmL6AyXb8JAmAAS8/D9emcmFIklmEU
DdRige2xd/VsjXDAhW+AIKmT5df+I/a3RHE7BJgZqoQcrnvxyE+U1XpXL534hlya
o5RCsRLVudB1lWwSXwT63W2eHaxpdwwTe8lgW/XxfvIIFOq0JiPxBpLyfyvxkU/0
fiMLyfCawUB5xtV1LmLdxpxyY5FrVMrXp9eU7kTbIJ8/0jF0FYUbCwWweQwuYcBX
GtLX/5Gdj17ewjpxXvSz2imGL6Oy5BEa7PUSCjlL/5GHA6KHl/IyJdNmLfhNcGmu
qlYpNyv31vipsELvFvI1KNL+Vybw3oRQ4zpCoHoHluB+Jpk62rcGrF8qsUPetmrI
DknxP2krn8oxWfzatT7Zm1xQ9S8210bvx5WGVVQN7bvnvFD2PZi7GC4TsSX6h0PF
Ub2EoUiUFS4xam0BN2paUxTYiqzjD73GAPV86xTXjNor8oZOm/mAtSvOcWGtDtID
uwLdmsfypSJ6ypls+xDp4XalVf+4Sk/xQiJpdP/6Aw8wAvVSsRe5G1sBuCTNp11M
LEbzEa3YpRAo4+pO+xiE8EW932h8fwYoOL1zl4kTV9Wov9Jd9IyrdDJKc2Yy0AbJ
Ewdmk/fEmVyPZSgbsuoNW7xrAWWZRv1ofdp/6/cIWtDk1f80R61Uuyi6ixd7dJ+x
OwZr5MuzV34rN8zPXYP+pKCIsSCWCB+wDsKD9pYTvRAcWVeimEb6d9+8G3xOdQMB
qx+1B9RWDxotj7t9wweHMj9yWUIW5Od07GIQPOJ7g2W1um8Ir0QSbbYMiE0CPqZP
XylJy+WHx9e8RgQB19nxwEVrq87kirGi6YFmbWlhbJHURB5yncOn4hXJpEc0VLL7
2DGGCDu32Q+c2qZIJ2CBRG5GJJd8IKc/1ztBk53J6kG856EH8ut4W8sJ+5VVHLxz
hAE37Cp06nfGRJQW7M97n11s7udrFfMJdJhSSKUgSPDBhtVbyqYekqVD25GwT1c/
8vEnVupEpSvT4S+n9PchUlXLBAoWGsoWbh07E7oCicM7FR77lUYfzj7OA+Yzp0sW
WWbAgyy2vOVas+RxvdnhJ3jzMY1eKPU46fJyQfSYrMpOtv1MIjsFIAu0aXRXvssc
Z8zOQhYbWgKiSWipLXccjmSe9EWWznW3L/eST7I9euoAJWkJ3AHowmnAuYxO7UUJ
XAPsE+OjUmxCRBUuv9bhD0Mx6EhpV80pyc2/owIsTEs7UwIWDxURmt4Y4GqVQZaY
wrK8GCR6NI2wdYywzvV6cYgLnj7HEzsAmcQT3RP+sFqrv0YNkJXpYTWO9v18+BKe
6Jay1yJxdy00bZ/Qgomb7TQAqO8XO9BS5zKZmCaZUUsngETqSt91Yi/0AhwSGAwD
pFzIwt3B7/oLKmgxIxAiIhfAN6LA9/00ySvFs2+Jep+U+eBlMoF2tdtY2mSKoRI9
MDw8pVx61tjfq9FVpgwwK7cJCxb6n6sn+3Nk9MVWuGgnMQehIademZ/MpA0q+fL/
S4W9X6BdzB1vDuSWipVRmYVS114i/AHMi0MPKCwaYripEBuLj+xhjw9qZmh0EGYT
lv/ZP6Uar1u36BHm1h4ygcub/wwYEH4Ci7qbPtnNreKZOFIc83S3L5958aA6wV4v
x5HAb5BYyGt8uKseGSXJQsJrdQZLsfbutHrG9r4DJ14OjO+jiuEXXNq6Ht86Na/V
P/GHhe/NFPZ+Fzy3V2t3b9lLJDAPEsmcfM7MHA+z9vH3a/PTzgFj6nxaYwz+osbN
sbUqJnpvNnm92czwt5T9o4oi7Si8msGM4NTXAXDjOxsB2qBjoD+DY/3UqbFKUHKr
HwnGzjMi59GiGQzQHxNS95mUXDqn6onJJf9Dkfz77dBIS+bMscdXt7/gd1Ldffmi
dyAyBEThpvSgbsYH2P/5u89kKLeyQ+kAp+YPBj1WMJGFcAjwBq4ICyKrSvfQm9JJ
QM2B4NZTzI5ubcxC5Gtt5KeSGWu4TAzumKavBRhCXSAzjACDCRGZSIn4Rssywoan
mo+NTBVHOLIk0yLT/W+OcAUw47bZBwkf3WNwKg572ALCmc9+Q7Wx0Jrlq5UM5qVK
Fe66BaWhp4mjzubsXT1G1aUw+4kf8B0V5bLo8aLEXdw2WrB0kB885fKi8QSLVfxz
KG462ukV9DRghtvtYbWtLK8LQBJW6Lyb1txuD7/RsPAZ8yuWTH/PAsYYWubJmqyW
StVtVcNUohnUbF1jg1s+9/2YXzgs4icR2g8D3U6p/nc9RjPF+QSHvZLfDunEwcIu
7H4P9SPV4nNCKu4Ju6PAXafHmrPMJJn0UIBx8LL2xe7N3SvB4KstPPLpOl1n4YkI
24mipZV6UdnebwUJ2VGUexH9MW4iR+s1RbmHqaaldtlStn6fY6m4BcPjLfS3X/Lk
j7+at9yZ17RhxaOobmlNAjD7fR1SRbBKNvma5/V8nUiBhUj6diQyXMNprjL98mnp
0R9LAcX9TxlvvR87l67/CfIhGvercnu3CrL13cCcVhlmLC45Dumm0nF+VINgaaBd
NOHmBHGqPk3P608ThfCcAVg9cmwegaW7Xm5Rqz+8b1XbdWLVsR30/XoAMR0Yr0tj
fo5gBz+d/PPl9Bc8VMg6qYAxhZh195ZBc2k5IYTU78DjN7yYKm1AbzGXCGR2srMd
MVbgwFFYLEInu7dUvCQ1OgPl7o9yd9/HwF6C1O/iIUlOK5tfzoUCXOkS9KUZBjZj
smwazgLRIc19ZbEhYCSfWE6SWIm4QyzPm2HAHbb3qcAG4sAWsnez0v/o3VnR7R9X
JjUx4vJTtBtTdTSyBMCVxu6jkTTKbMY1bpx84M32CIt/1OP1AHMzGgtpw7V9anym
G8LgElnq99xSVzkofw/4oWFY+azgOl1KaRzBx3EK5BmyhX3h4JcTi0tZZ+sJwmVx
ajuRmaL73PEDu535Am0FJhygd2g6S5Ziv/MiejTYb5VNhGnlNLLU3mc7gzAf7dgB
SBpuIwibAvzsOzKz8tlkwkU+ULhYhpzE8sfkoEtJ7usVAzF/HBrrrnYzNYS6DqSB
lvyFCz+i3XK4LU7UvDx7UTaPr2ZOYQznq45qnlPJbNHsJhOIjrI1Mvj1h+Vc4O7C
2BVjHISei1KpCWV8kpZDwvvFReFIuJwTCCuGy8+7mBXMJQRsxH2ErOIIStrHSHt7
9vmN13YMiyRXcbTji9dnTSmVSXVF/RVUjnU5LyOBW5YWwaqXMPHrITG/B29OMeEc
7m2rGQAf3xDKghe/rLC8wjVLfqEbqeoatO1M3NnSkp5LXzf7BHCrK/RLqQ0wrqpg
aDS59iZAOr5qjC4LC72qZMtq2s9IdZ4KkmejQ4rn+82YX/IBJeTYT6YlwdCxJJZR
sDhWHKMECVlt3iELtfncW+S6n3AFYCAjZFCKZuMzYy7+hknMnV4H7/rfeoxUvl3X
fXGRioKfv15yWFfGvKVEIsYppfQ/9HZ7IsltSo1p0Fl7+uy3XnhqEBsoEqWXDoPR
ZXGTJtg9pF3q/byBZpKT76WlfYG/SUoljbndJzfzq1BxCCWGWl0Kl5xLhZEqO+ZC
9W69iWKaHQtsnOC63HZ2P4BrvF3KtZ4GXJXCRd7ltYqWaZqMdbuUH5VQDD2v2JU4
c+weEOE57ozFSbiA2uzn0hqXSSPu+TOPTpxIlC0Dmc77022E18qL23eXt2+zotos
0vZeEAltxJl7w5CWLSlgqcz4oWgqNUxa9IDQK7bjHdxo+EugCgji09mFzkS/Otbv
FhJsN84HWU3Dia3o7o1izEW2cLd+G6yRqX0o31efr8H3ZzWKG37yk72qOqgEQb7t
Sc+f1EWgbqO7KGkSaZrHFDNPUotC0fTN5rVKCGtm8EK2IkMmPNZL9wCD7hnxlz9U
L0PSSGY4eIbs2sSsikBF5VnWQa7up0u3TDCMxZYJa2MLdifmxWLLJ3sE7+EmWrHf
WXBgFAwhmVDgZvKSik8fmY+7YtqRRMBzALamZm/rdwcft8HeFEJ1QV9o0NIs0IpE
pMlWPBymEtViktSHaoqDULTkhFue+aXYr1zb/ktVci2eYi+sVm4AteQcZgoMnVBx
gzQpX/dqKe0cBb/Af7Zdc16LiK7l3TBaJ2/+EWfPkTDGco5Z1Vl8Iio1+3K5abdr
dpSSBQC/MHXEQSrsALY8rSLRwY7ZL3qjgKtS92NhPHkZBqLCwJEYDGchj6H7vl5m
xIS4POEUAQ0I+HgQzy1FFmTxpKwfMpXYZekbvxtTMSRHTketPOpt+ZWz5Z0VBcal
uREsS+SrPpQP51JM9tonbC7edXZg18Mf10cQcZJyUTEa5UVrgXYczyVtCECbxGCp
2upyVJ8wnLrUSLECU7YS+yaLsXifTa1vyD4bKUVSrY5g9p3Yj8g+I+EnVzh0ZOKH
70Gj4aoqAvG+yKqCwN1agcC+MGfvNssJplh5jRfzAF2n/aa5Z4wf6IEAHdTfRtrC
Hrfh6dBXszVxz/gwnPY38KwfHu346HdV79scD5H43x/5dMqKo313WHGf6+DxlWKq
YSxdnSwO9ssgs0u26h/iMyEoiEjSs5kykqSgsz2aYoFJIxjWS8ZixoXO3fMPChB2
DRNnZGdzRyJ31+BzJekO1ewKg/+zJzJGMrgm5KQuz2NFHyXek6ZCtVAcPus+yC3O
rmGgBo9IXPr8b/loMSuLhQVTzxeC90JoiOJ7TtZ5P5pflwL1oYt+eVwirDGnEmhB
PNhKbXYkZG6eqzFLys3HymVJr8+ASUBaCgb+9RLMDnguDgE9B0K8Y4yuOG11oTtQ
sYyoCMqDj+TiAtChymxKYabItc0qzTDkqyjbRc1XQMjAzRsU5auGfOpypldAmpla
vSFRmzoUS1m0fs0+GhONfyKjduSWFFdNWhnNH5mFxI7A7J5/htGKwdLbyP6QqJ0p
DlaOaVwl/0JgkYOpQYpLXjYQ2oHSnTP/o0o3EUyuIUK5HH6gQqRasX5fJeqN3wMc
ycCDxPsEKJFkcRNv7gRswFKDNVUMr0D+2Noa2ZiDKmf43SfJQMIZY9mODvF1eqYg
D4gO2q9PEIji6srZpaQPqSRldQtkDt3xd47nQACjgCHQtE0ZXYEzHgsJVJwWDt3E
cob3bQaoqF9J6VS+KKCqUn2vuUB8tmaayk6trylJh1NZYTFTVmVciRJYcK3Hmirz
IUyvHBfzCXf/54MzVFg4KTPEQlcAbittWngH5EPctv+9IDLwXTIGxqYI+m5QhVUB
jsdUD8kQA4qbmKXgeEZFAbAJxEJEGw2je/K8hwmuWSoZab8FA6SGULHzeXmHW76J
rska/dEEys8PVX6pSFey3+G7UDXN8WP4mkcYT/m99yOrcWwmgadBuvOZXEwP0hCo
AsCX1Rm6iWIEi8WgaTR99mGmI6OA1YDIl/rLdCGNxAXBxdOy9t8Zyh6bE9n509Jx
tnVlT+SsQU73pYW/3qEpzTebTHWSuhCqsCrkR32XvRI0wA1i9ATNOy1apw7P6Bq1
C025bAGuxG2G7DXfbu17P2t42CAxxdPNkIq8s3qVHeUCsoEZkH+TVozjFZGZ7ezW
fKzrcshpz8LwF4ktIsO4ljkFVXKG1q1I2L2WengTimyiM9EI8WFSAXn+80QE8FSA
wDtEZWCxiB850j60tK7St2uJ0FVTb+GIrm/tkD5LCIPFV8ifI93sURLe4qmmm1qb
V9yNoXbA/1qvnlljX78bwk/beGzHRRIL2h2fZ11ByOiwwn7mgPeUOZK+6+hainlP
PbR1MLDCuFFiVTgqLabpm+a64sJq4JUmDO5ddKgloyE6JyUoKgyVJbY1/nrJJ+7K
gux8RNzSrLpeDgcslg9J4dEGDxEueSIxOtoY8QEnbCiGbXcV0lo7onsrt25wNpka
CwkWtzQv447Nit9QU+ajP012QG+GcsvRW/1pJ8z/ue8Aqhk7hwlGvijqIn7Lkxwj
sNPou8HqxT5x26a3KDWW12aVCxF8IEQUC8wXU5DR1KpoMrujZyKUd1rZMMi22p8Z
4OHvy4IYcUeKx4fQiwpPrWhmGtNVtMgfezIH7TKY8pV2eTRyKvCqDhWyZUw4wtul
Ka7jiIW2jUO0f7KhcY2jpAbM9Y+kiKLfmTMaOHnM0H+5VkHV9urU3jFYxKEcNc/R
7X4PJjtYYW0jjP7iGsfOqUMh6wMgTcAL7WzMzHIeAxSNpqPuyvXrTA4GBmBJhMJE
4cA74LvMaanFoEIHNLqzbe0A22RG4auj2REH6UM+ZFpPrumTY0p+VYl/XvfV7CiJ
BQoRvQSNyERXIeBF8gE4nnTxSr8IUoisaBoC/IrI11rbIAL0x7RmK93JZ+dVFgeU
GWnVwGJxFCDIopHXLyoArFnXmJqJMgiZIrGEQtFbbX7fhJsPqFgjbAmYix8sIwvM
kEeTYW0dAHcBk9h5lMiizVVzhAV6Lg/zcguu7uSjUpILZSebhVRs9v9POjC736iP
Jv957dxC1ugpPHRpbzpMT9j5buHD5UKbbUDWFzLf00HNafinzbdrpxCmnlPJWUAV
YUVPluEuanqMU4IAPSvJ40OZs6d16RVUGmzOZqF7oSuDFznO6h+W+ATHEcJHLBR3
hK+zlvUCNsE4HeXPVPNkwD3zfH5g4n8AJ9J2f61PDHr/Z0mUiRzDMgYO5DHqB4qm
XakPqkLDKD6czCWbLl3WH6lKexqhYe9l+U1Baqf3yz2u8CzisFn8LLenyJjzsekQ
RVqCVRMKvJwSj3H7QPnue2kc+W/LvIJlx07uogQTrVklY3+RPLkq5A7gXa22Q0w5
Jc8f3kIbOFkPg0oi51BSRRHIwivIHCp/ui6+VBI4qRwoZFUPnKOEmxw0moOFS1kL
lqBqR5eR3zywrmzlmqbqRDFr5+mShN3R8FsUW+0ExzLTgH2hRBlXV3MkYp27x7FX
+/GeNbHKmuusFlqLw8S75GbkIj9eEt2xlrXg931feealZUVQTsk1NPNBKASdq2SR
nMZG+Xs7RkIN2u6Sg7glBaOiir5RphhU7L4ujgWRT9Q+DOu3ugWBpF9acw1V0FRJ
SSWBOyJjC1HR53x9hMAzw7XpIcPXT2x2bNuZSh9SAFremxOF6ilShcpDobFh0/eq
kFSCNCAjh9f1kNoMuucHpsDtIYe2fYFyJNceul9o8GFFpWgGyGqsb3J5f24KoDhH
iFCHXwP0VRzn6KemfV/w0AuAxpike3sFsJYVSaEpu2ej36F4DlERDiedcMCYkGP/
IE7QzSobUF3yEF4xd7Gp1GQWz96ZIfPDQcuhPCELdFf0y5V0BWPY60ie28wKz477
sVHeFZmfjucTeqrOiRFWnDbldba64j5X61TEoMwSW/aTp0ISTNzUiyP0QZbMyDem
71FyfrTr6017xbUkyt74rl7znLgOeyA771zH10BlUXEofyXq3m0i/lX7JoaXUcOH
eP2IqV3ZjWYQMuocHRPkiKoOxu58R0EV5A8BlBDQsrgQ5hYXRlmpZuHS6BS+nmW5
5WHYaFmCG4XM3R0SQ09PZcFKfQokH2rrPOUG2MivVetn85Lwum4vs4z5wqMcjZeO
4PJcuVzoUO6A/ad1hDAy/hjxN+SeYAlIdFdEYsWZcPmfE3wr25JCYXa2XjrMc/BB
oHq+4QWCOAOnhqhA5w/k9NKovuq1qvflmd/V+IDbZQ9Yaas36+avD7AnsNyVVYsv
5dW+k/JD6rS8sJkhKjkByZzPYDmgfhYSKdhKR6qLTABbx/76MowrpoZ2aLnYTMQ3
+Gei+B7FiHuvuTLqytVbPRKTzOHdqnev7tELTw0km91Wi3TZpHgjqIfzLPapAEkh
jIj4SnevwkG5qHQxLv6EhbrwOtuqGIQyoLKzmfI5LhQCVDNzrK/x9LCPogaBI1MA
exu7gupLeOtAwzJeqd5/MoaltLI2js9022SX2Eq3uGlLbJJEo1wmoyx9N2/giozl
st81HzUkCe6nH2P+p5A9mHctsmvj7yCTjWonfTjk8dOl6FTuWD7bo879Yq0H0hrQ
RDRAj/ZWkmATx96mwVvLNV3vu6PH6Ya+8CWKNYOEm0JU04cjoYC4cVcj2AhWeWQP
H1rgXh7C23YtvEuX2TjiTagbNVOJIvH2dF3wYv/b2Ob3thEgXssXXo0+mK2Earmw
LMpTyUFXQ59owtwSH3R7GEotqIHBG8Te1kCjRS41ArMfODm5z4tSCDTxcS2jIf7m
fi3iEDmZSRbax0p+tUvF5TI/gTKd08fGt+66UdcLZGIbb16DG1eplBtQqt6yuGqV
J42yjiJfkUMGR5LLFm4S02r0P+bYEWh7Q/rb8wVpiXbz5/xdJI1R7oCanoIN5mZz
/GkeaXmRjWf8ImebuTYPb8KlAp4euLkLHdna3meNGwd1q8az2aH8R90BY+jOR2KI
zJr4CnDtovOkpGkyKRKpQCu2zgv2mZES/UYixV2zuQwqhJ26xV1M0xGoKkqqLArR
APNkdmy+H+tDsiaPXd2pKQgecFT3CtlQiI2Tw9nQbUpebhXLUcDLOQaLYT/UxvJF
hAFlS8nshF9yOr791rILNGl0rkRV5aavZeKJRK2k+mEERmcMI7afwfQOO0N/Hqao
2a/IodBCK2M2N0bLmzhq/8qVkD18P0noBpwKrbtwWeCT5wKZZ7WkNoTSTboMIjQT
4PSkoShrTsoVjqO1TLmQmA91Jmly5jH3ARyJeG7SfvDQJsvV1kXDvbxFZbKrYdqF
vtggX5grG8dDGbNNj2HQBxgsWFZEoClnKbuTwCYT0UOWfxTR4M6MmrCiu/74uvqE
0k0wiKlcC9GvrqEOcZL9CJXOEnkfHQpW4I49JQjZyoUh+E4gwLCJW1s6XdUz4Y1u
MFAk0LkU/vxL5E808HZtmWnodxQcOvA5PNxk3qpO8xk3YYFWV8RfwytGe2wIL16g
LM29/ineaXb0WR0tkyvEN4raDijxhVUCaJZEsnI4ip2ZRSm7F/lyiilnqP3bxDcV
AmBAPDNr1IOvshstef2DEm72A4gJvnLBsBjA8uA+cH3ekd759q9jJk6urxeVjzZJ
BpD3A2WeSrHY9k7zgcATAQODERuz2OTEvxl4BqnuYffmTpgWqwKXOZAv9gP0dEAl
awmiutAdNAYKYM8ookj3Mzj4jpwGgvvb9HemP+ODQL9VPyf7d+mDqb1zqxc4W1L2
whaMeMZsh/GsX0YAfkjwM6R+/nMGvKWxKvRXiEjTCiqmjnFrz0JEC3m1GzW0CLH6
kfdFU45QBL/7NhiPNNeWHhYDBeTHbWLCyt5EEUumjIhfsjmTtdBEyZv7VGNNzjET
ZEqRIq3j7bnDD+SlxXfcJwrku61DX+jfwNlOM493cijH1Uze65OblEFr6TsQDEft
F0VpVmvnMjEm21jd4RBuOok/uWRznfDJDMw4jNAPcFnD2Qm2A1OH43xpPwCH+Kxr
gGEQ7qZyIchoqU3URSloHBGlPzJsA3VZT/wzrCm7fLbiQycOGm1h5zf0CJ6xfLYV
P40jxVCfuo+h3EVY99A6fb4coUJshm3v+OoF9OUWdb714VtwYWOZs209tj8qBJ+m
N+gMdC44b5H9gJ9FasEYL2lUm+vk29gAq96qwrtXg4eczCULVGLm3VthykSfE76c
rs5LYcIgqUE2XtXsQHIa20h1eB6I24ej2deX5km2DkOYMYHiWw/FPyAHwSdEjSOx
jF1JCexpEFXjdHBLLZ8q0M5N1DtNQlv+Ax39gNH2rSWDKOcdl2WcE3g/4MuFFQNg
KZE7s572SCctw65OFsO37BokNP2zKGdunoFSNPkvKMsFHSxk6TRxIn7cgWYkDwN1
e6suDRktNHxgqwcy7GOauaDuXfFa6ZmChZlfhRbqWb1DEF4JuU4/MVGV1LTDv6rp
skc9hIXnrD4VNouD2Keh0nYQUXsJMtCFhHriNf6JcpsbQFaivPgFMfzb6n1Ld5ha
aa5aMz7RJE0QsQdbS3yZTl9DrfAo9/s/XsTPnyIhVVpDz7Z2ccuuT6hsK0xvMhhx
oFevbOZGPDsdDXHOQ44BxQNh19bn6BTGgGhdCpF4YI0yr6YnoBRHCg+HpeECxpIy
AIxeoG9juMgGwICKNdCOJn6cYDMwmisqW19q/W9FSIQZIP47mjLHZxqdg61WaDA+
oQZgrmH50p7tIz4nXWBRZZkUXNXEiWIO1hlj2ozVHoA9lnDrSrd96ovtIYQJIoDQ
SuRI2q5iHjnYZslk6obFM/oDgf+svHFvjhu1TsFGW970ZhMP5bljNY0d0aJIvxVf
8T9hrxAoCCmxM7P1mJ1/CQoPCNArwToSew7nTX0x6HgwCrCInXM/xv6kxqUyKvhg
+M2Pa2nNHpABOvmkQXc8nVVN/Mqg18mXJocmPbMQg8N44geoWthP+DcLX7mTsFJN
cx2XMZVrc4wTNA2r7KGLWcoV8+SKMP8YGruz+kH/WJjOmAO2F+0lrP59n/PquQS+
P9/4EVqKdf5NqyNi08kvJJArc1wWlFKaFbGRVPiSsPK4h1wUrNqbSi3oDxMCBV4N
1sfFNM1aw39+kfE233ciG39Fq8HdcAO09ZPFWFNFIKMEgDhmEhmsVgSgsMcjcqip
UsBoshr8GYFp6W4a5+nhycJcNpWB7KbLeRHMwBeSiNKnIayhc5N+l6+ssN0QWmLy
7zivMJTN/546+hER6Ljv2N1IIARcbpRMI2qpX6MEsKJvar5VymxHxbMfExEgmmaL
kJVUL8GOpPmgkIS4m5cIKSVI44y13wTtpRwhjx01O/xc9vZ1TLkcpWrjMNXzqAFB
wx2sdHFFXoJqJFfOwyxCxNEb4tNAhDSoAtZfWqfRlTnBO7hqx7xqVRfXycFatFMW
R0rasXVjF+tO3BFPqBcSUwWj+Gbht5dA70meFqN5SHt3VLPAByagt4ef8ywGcnSe
p7Yf8EPVCFgCk7ft6ruozpKfo/lszDfCqbkbFaZa0/ikYJNkKNaxPdZYdohkfdPI
r24Q65CHilrxMT8zDyujcgpi+CFHUpyLfCeZy/bjW3uTJu9wcmuzD/ma+4St40a1
enoF4b1qMBDvkX2Q0SRHi+zA6f8/bEWMiPF7toZjSFimsGUow9inTSIL75SlaDGH
vX/YBSn/4Q9PCDoMrFmbJoBlLKkM5aZ4ivI35laEzf58tWd49ln463juO9FtNemA
Yk3kGsoeuunPDVivhHzHG6Dd90Xf8qmPFOSU0+yrpdNztYbolAfYvfDI8OgTVyG9
HqFGHbuO4BlJe17LoZcByy+Zf0LsDegySSNAeUBVxQ49pwqWyUhG7JNIM5qBGHcW
AHSE/gtqqVqCNwk3TlW7nIXwfBNkm/9XGris4cOiRAy6zcQrogVyqWcLHP3avo9G
zU5WdW6vaC3l+b2Uk/3HXALA4Nh10wUdd2s96eTgzw0/Cfw1kq5J4I+aVfP7bSsT
iApq1gsGYgu6lB4GOygMyRW3+HQ1mbqBhk0RVlDXO9CGCJ0jC86esbXbzWzbVH6E
/vzpNuSP1jzygTctZ0eXFEfraIgEeFTM0iNmu3OwAlUIHuvLcoqHLv3xCwv8jRK0
ZiZ2nNfJA8seLyNX2vAYcU4ppy4tVhCGP6jTWmi4cjnbDVUJvJwnjQGWzv1FgJPf
SOLx93AJ2Js6gLvY8Rq0Dr1hDcAgkQPVlBW9YPOex1RAmg9hdkdvhxPdm+puWmvn
AJmA07j8HV0CeY0ddEEziv4OR3dOVAZNb7PGs2DOeGe5KV1bCVZBByU3QOKyfzge
TjNwFp6tmPeTN2n4A09gXk4+ctJN1jUirQJMormUJo+38ECJIKn8O8JO8xQ5hKGQ
LyxNl+XIXzOidvYuQVzwtbD92w0hOSwzwvsxwp1bCOl01+n95GdLgNmVZW2vihsK
LCVAKfYLld1yiXxcKZmmtkSGTFmfIwNM3tEVo2o4WRaHrV9z/M4S70xYePo7gG3B
gYvOx+5kPseGqkTFiOVNo6WKA6hnlLGXJQGEnsf7zM4ZwO3HgmyIqeiJR2s6Zuxn
tCeKo8CsBudi+7UklWBCO82F9MwkRhqX4mWAI816Cu5WoDJmxPS0A8W5gZ9+8h7B
AQMyr9VvLnCUS8j+o8L84Y5LH60fFcpx36FCn/bubKS/E3Z+6jYwCB6SnLszFULk
25A4EUk593orGx9cgWJ8eYmEKbVzmXV+M1UTglxTlXL/q3CgUO1LzQktpCq2av1O
5UrM8etYuoCPU5wEYcpK8k2KmjmYIDKWFyHK6PB2lyPGnjkiRDnb2/p29Lx7PaPM
vpO0GSN5/Pv2QPGb54k1EyeEq4Qpc0r6LR0N+H9UIGC0eNmBKuYW6XswMI+O41Ph
CXlcO0u1ctz+nsPPIYucRVfGTsFOL4O0ygDQKi4XxbMZ8sUtz3wOY55QvaW5cv7L
nWn0BA+6M2ryYVEKH3YsmKhnsdYvZgdrr4ljuhjYTXKq+CVj2HoYvjCfcbV+IRQ4
bOl8HnYDou4uq5AaGcqZ0tUlSgvHZK7l1jU975wxRTycfhjowfjE6crr1TFfJ961
1t6maUEc1ycQGSa0uBZgrwl/uIj/StoMHl9BNvCvd086dR04o67DQazxV/seEaAf
lVSeeNU+OfmK1JJdQz+Qg842+ufu0idIlLtppLQ6U3dMtWn1QTFOLcpLF5DRvMc2
mV9eD2I+f9JYtuPisqEve9RHt0TVkzBY9B+buStC4Ep5SKELNajesM6Akv8m7vfU
FIXSbzdKUGRi1VGsyB3zxwT55F+0s/45ZI2ymQdxH73GIraUGXO9ieYm6rakBVcs
3w5DKJ0mcTdimi89E3D43dp+W8Y1Zh9dtw1KCYIErQnu9YTP9dckBZXnKKkFMZcr
0lZYUPOIwjeka7F3GsBMcmEFDEhE4kG4C/ukxU9hkQDTLtGx4wAXq/tQkfygmgf9
VTXfuY6GnYyuMi4yRoUzaswNARGr03nEqAjlv7hfAwkGxKs/F5DhLxHdQFu1JqjG
Z6Uo9w/15j6tP9okKiWISXv90gbUzyNaP+w9UAvzZv4zTkObpcXaPGFrF4aj/cOU
cW6cxA/lqCGdKfF/2MyQh0mPeq1GoIke8JGw25usuz6Mb4tE9jTh0aPUnjkIv6zl
RFr4xRfNVa5EgSORkWHHy2+jRbriCpazADWpmzDG0LvTaPRXFD4NXIWFOKdiG02r
LCXV/ei3NDM9OrE0jhrnAWF1Vy0LbmXcV4M+9Mh23uBd/Qw2NBT24Q5zsQHMmTUn
7VflCy0XukgYigTx5R2cQ19AZdHdcrYPvqlj8DqY/cTJeDPtfj0P4U1S3yH9WgX9
f1EbXe1Evbpb3la59Ti0bAbWvOhR2kQ30I72uxQ1Y0pqSuamFDTKeDQC7xwZat5J
Je3pEougNDL3RQGb6DCC99mYDK4qWLJMV6gE/rbgJuLcxYY3INGT0iJlSdM3kGfO
bbeBpHtk/r5r1qvqVA9PY5VkVjxdBfmLv8IYwnz/MDbAklxwpOTeuWmqigxvAbTQ
hagn6V+t/xJVJRO2BJxArGJO4jsMM7Adjgx3fNE/dwmD6t+8EQ3nWYRVd4+aa4ze
rCr22df/xF6+xsSzmpDRn4R/rOjF2xJkymxjhpfE6BjG+Pwh7LqCnJF1dvyOFY4r
RgUwPNdIOO3nILhYuhTwVaODWzUSbW5uXTQeffXxQUb2hVX9wC3U0TuVl5sZ07xg
+JrmsJWV0GkSqgrumXoItuRuoikAPBGnrVxPa/xBvLE2f5kRSVX4SXPg9ZZDSL+x
RweRyfVeH8nEmPSr0qazb7L0ZPi5abXUftL6lseFEUKVQHkzdyXLVlRb8f3FO9qb
nQQaRlyHaWVW7uT5j2Kyz9dfrV0lUbNfqIJgTvH/5awagIQkVUFl/G4c1S9wFqJU
QtnyBOWOOd6ZOMbAZY1uc3oAmsUjuBjJqfPQc0vRMofXoY0iz+DB8cLrqd7cDPhP
S9ZY2/wbCuU0IGF/tbfDVyaDFfb+2Wt1fPfT+dG1TwsSmrf1br2XxRi3kPp8lgNW
6or2E0/HpYzzVJzVoppahOJfPRgePr6QGNS/+Ev+a2o9RXFeDnbIoNOjCdEK+lbV
itB2RHogbOrqJ7nF5W53s99EAPxdTdQa5Y6UvCAQvci+7KM/roQzzdI2KGL0D/0k
sbwkOVWRWhakC17IPjux6ZJ3FdZdzpNBgdiPla6iu8M/9jdaUWR6XAPvElqcc2Kz
F0zQWL4LqnsqBI4LqoICPn/QIBy9/rLQOxn7OSDn+kmAjq+Ts5jAZNLqYdqNBqE8
G+285+t5aEKI6mc0itKk3gk+2t1skHx40V6hUwSxGhz55tC3Ggsgdb2aUXlFzHdq
8j1/5vW4Uh8GFZ70EJzQQLqEO7KUJVFuJxGRfWBDSqcCuL0309+Qmy4S6MYVGrtP
/YrLJQKg3r0tDnTvj8Wh8/8g73kVMWCpeWoGLdmlR7pswIymzyMCxqKuFx37CWyH
5+tBkmxHpHa6kOWRUFva2L4HIywnidpxCefZOTB/21LDZrvH4yc94SJ5llMxYtxK
hpwfeJeiDerY5nDdDNGZmdsw07vvRni8QvN4UeQvQDKDTNgzwF86pzWqxCSG7kIL
wHaPwMN/SnwJ8fsK6qM6WBTGCBxTazBewtWrupvX4AZkzL6F5UT1L6rtDuLg93Iy
wiAeNFU0IShT0S/UNPuLCnbDdX30Nm3c9jPDUWXEMFDi47j8GIU+fA/GF4hoZNKX
ZuZdkzmAdxwaGFxuy8vbFWXWHIXl/D6lcRaG+QFMAHBx1lB8jJJNTxlN+ISmwp7+
EeOT0WXKDe2XW7HF1I110HMELlyt5mgqY/wSgWFSxe8f4tXISlksd9x6T+KsYtaC
S+UkvEkixGM9DlAqxIt0hu4vzQYH/ub0+stV1tH97LC0cn3U1PYZ6nJ7cICNw60t
3hVf+lp6MIgPI0LzIM+FssSlMMGtF7c7g5wayvBk1TyEkLk2KRxp4Sl2gAQxTy92
qD0KkOX34EB8ALzQhNnsgLV2ygzW11NAE6c6WYKF8cEnxtVXLr2vLH4kXsgCHzGS
IUBfHTE/afnKZapYJYlbmdYr61uOJhYKBSUtrAgla8sG1Ltspu4DbpJZmB1flAoo
l8eJSKbibmVgnPJTO/eJYktQEWX/cZdoli0Oa3Y8ph0iBk2DPlKnUdLf5/VEMuD9
hCtsEHuM9MTaPeKAUBX/c/VH248ROgfPdxyv/kLAlMyzbiJ9XEq1UJPPCWmyZvti
uXkRd8kzICX6kbvvZEnwEAXAZtV/sBWUJ/4xyz6tll+daAGkyzWyerLtG7jb4fne
H2X5JhjKxn2+etfyyejoKKMBoTLbrBn3tskItkZvCl5oLAaEmObDRrrmmOsSS5Su
+sqMURBm1+aA2FMkBQGz/dD2NxQmw9S2Ze+M1OsFUiF87VTaUeJZjkQDmxfSL5pO
8wySG/SWRmUXBDx2YEB7O4BsYKHACImy9d695rAU5SpLGCwwy7SfTnuqIPkhOFKh
Vtuxwe0dnJubFvISu1or3VsOy+XrWRq2VK9D42yy80RmO6HA9I4rto1bfQF5TMZ9
24qWBjqEEE/quIstO/3Elaa5MF8bvikJJLKqitcun50hDUE8GEyjWkUVh3ovzwp0
QBXSVbeTm+dEB7ZeSaoNK88IUjdtBH5QIHgGkdzBu/475SzSEGeqkaRTq+Y74/FR
Mygas5y5ktdfPuMoXZ4XYLhCNENCYfrzV7As7vv+8mC0ztfQYcdYv+az4sdp7nrp
5ecX7xf4ChesjAGkq/C0HUoYa7HvPyGg1PyLuRk2QOPa0EL0B6bYFHHIfYgMivnj
ui55sbj4BLkaxHurlvigEtDVbFR69kOOt/dzlQUQTWZwKSWRU3k/PbsjhDSAq7rG
Wyi5/iAuegeU4fG1QABYNznKOcJIbs0GUXMbBerXHI8odMu0BWvuPrsoF70cD/4I
XggGL4Trc84CAKDLiQa87onohYSs9mhuvSeNctAhIPWhoZ9VPipT1M0AWl64H6mR
DAyuqQkougY860GvQ8u8GVaeFHGO8PzCzxYpkKVfU+Mh6Egw0OQqgW7deeCLNJio
JKOQV+uXpSe8VN1FJWaQ4DSx6402E3v2cbN4LKScIDY8CqXIly2Qz9QlXyKTO2Bm
Pc7V+rPOxOA9RyhmAgrp+Mtde2l1OnNI7aOudXuPX31tbGN/Ww6b7VTgYzJCueHQ
NRLIGR+rrGGL9Q2zcwH4Ib7KAbr5MWvET8zjO987pRkHUFEA7J9lkegVKGILJhv5
B65EUitdCmePcz5TVPv4Cbse4FrrmT/YuskKr5CgbICMJHs5OwdsgxwzHF6ssFub
qKQVLF4mas822ZyqyVYBnkpCa2Fzryz0PFStE78i0JWWjhtifEpOkaIE7CppBek5
iN+tcVBMVj08ctOV58f3Kpd1vM1KQPB7348x7wWhQ/4uTn3KvSnOSHon7lOtY+BA
1nFXaRvDWPrejXE+j2kLM1MeLrc2C0lLEvpJBjsQUvjOUG9SRCmSRHWTxZ3J67Wq
mDu3p40GVejXETf49AnVWZ6OGg3uXs9ANpVBBsyTv67rtDUTYJBS0OOhTzPqwoG2
dIsCFe5qlm8PefnwXFLoXl4WvhfxpCkuw0Ux767W/YVNUpOeWX178LNJ/dbnaXaA
+0DXnLqYxyhyhSI+jLtxua1KGei7fe8oxrdwJj9TpuN8lhX1pe4Sk/7dAxv8gHrA
wBPsfaL/AsKednm7FVWal5CC6oZ9GoG4JlqGcxxzevvk0q+yhJL9I0kDggVFxLAb
wT4bS7khcB0AnzLMga62c6EHLhw12pUF/2Ps/xNPGirqOveIuz8VhYhgL/sCjPJc
cpgs/O1N0Tib95wr9aTbiBcPSUPYKf+bSNw6mZGfvKZSPwj3sPJVsYLEVRFj4nBg
ELQSO4pqIe5F2vWmLex2DpIoQssMjzHSFMwgVPmg6wDPck2TX5cUG7W8WaFXHg++
nCo3OF287iUEtao3cB+o3O/6tiEhLQRsVhXwARGIfa/xF1/lPPepBZio0YEs/XU8
dehMbXcLiH9f0tzq1uzvIEzCi2WhtPWlpIZrJCqnLN1kcsj78iJIDsEMoWxwvb9n
VQ/ki2oPQR1M8sbiImRJYm3xQi2aiis1W3skq5XjLQr9OAjA1H+hTUyAZD2Qmhom
dIkSv9PEbELmyUU6Yx19ociw8YY80Kv+L6DfF7kwP+zE+kDe/fTb/ikzwMbqveqn
UqoEN8H1RGmSZOSYBVQGAnn8QKHrWsTilKjJU3RtS0amFic3WjT6Gvxez0TtOwdI
pn8f7I3/i+vzc9S5+D4KZKmZ7lcJgs9E4J+G10N/dFVR2CYiLHNen2LGp5VyH8Xr
O+lT9a/Ekx5cIFEvtlbnDKFp+00h0j9E6eF+YxE4euRXdDfHUEcV8XFy7oqM2Olp
vENbQwWbIKbG4aSZL7YFtmCf0ZZKRf939SKE1zEhOA0sLKHuRuiIaxM+rH0DqvN4
6ZmGY0GRsTfQ10iXmqr5WjbE+85iQM+1mlSJYrXICngZ7VYWFvgULW4v+6+Wd81Z
vNd3V1UJC3qqm5lIIQbPyKSoyuUlDaEA7Xu+doee4cHQaJzKDnn7BMVViuu2YpvV
OXnMO3BpCKohpXlXN6m5lS5kXVTkaT2USkkMS6ZrzZvhZWAoOGOkzgukQZyJ3hFE
ek/+AGIyOsn4RAYP4S6jyhNwJ6H7FSWoHHjV8pNt75jexUN1MNXJdrj1uQUOkqYw
haBc7Z/bZDR+NvULY1W4ALu7jh9OR5mRQgXoYVr4ajsQRX9znwleEwJYKQXlT1ci
oibr/QiW+Rx3VTfYqB820Wl18ifVVMWswqSgOC01gM/FaHCldKG/21fIKNwSNFy0
YlNALAODyV7bK1vWzDN+LGBx7r8wQKIctr2MekY7zw9c+161FCj/hUHh4pjmSzfj
sBQ+vqJBW4AN2vDMkJGyMrfO4NSPYrqJ/qpmmUUfjVQBhFzcoqLXD6+UNnweGhDn
tK8OO9hKWugDocefmRWdCZQHzRqmSubL2P37AOanb3qCL//nHksv3dxYl6DS84h3
L9NPDpGsieoVkNaZnAbNykc6jkvIZu/m2yZq7MpD6KbkuN5EEQ57/YJSOS/K54Dn
rWieAHY8Om1Q2D5hm2f3nkokQ9svLYWe50gxSXHi+fMsgYqS1ckR6CbDIn6TOLyp
2fyP80xrmebtndkTnkl6hN6+TjY6ZlZsAO+/a72bqm1FWP88paF7xNf1d7nDotss
28HLIz1KKFKA0hFYLLXh5y2JwBwaQmHzj7iY9vFYYSJDl95f3EgnlLtQnnTjC4lS
4/AsT2dg6dokp8mrkX9GWJUyM4JR15Lf63JCDWig5tXaDnc0gTBtPImKNxbunJE5
QbXuiioGRgJWNWNVqyrJ4+1dinePB0XAVFyqh6zDCbC3Po5LG8RJ9dfUpT2kCaZq
20l8tO9iorm3/FTH+FcoqV9HrKWbeArMIfLfePrjBs21Ap/3tv3cDh063Xk5LjQr
EvvA/QNQ2FfrENuuPJO3rGBKDOAlcgbtbIwMeTEbFyaO6pCiw4bVwpA+kcKHLlOu
FEj1qdGobEcRp6jyXeXTB8El5gTuR9Ea/LKdC4rAeUGiShy5X96dbEWTkaMEg1u3
TUxkKQf4kGOEDeWe7qGdA+ebsnf3jsfjQnCpQhUzYdMMQxt9NtU47WrfSDk1o2ke
pzCjIvPGVF53DTCuJQnQ7F/MDVc3+pTd4BcIxu4pJaMdFcD3lOKZftaAt2bMbymt
p5Pyz3GQMmRunr/X9CXnU3nx+bxdz1s05TZs/b6TWmkjNL79SqLJYlmeYVYTI2fO
MRrfrZ/TCUsU+rdU6/Jd0PiFW0B0MT1nT96qRHWz1u5Xfj2gI6SgjGo+v2dX+SJq
CI1BKGtQSdNZ/v88p4ZieZbGm8Ju8JIiY6gOYIIDwrPMxhPs4i97F4UJGmJpQD4/
0ZktkhJL5w0xy4QsXoQyw35bVDWpZpizm3zdjWwnuwMVnrqNP4vcpPPOZdII1Uji
Ef+4cd6OUopgslzql3HRM4HBaO4nD1Ic6ZuBGrDA4A+okwe9HkRrzOS+xo/BxOPX
Ed63FBr86DR85s7d5MCXCtN8R+lCpHmWk6qYmu1QBtcJpTnY29imESG+BLeAr3l4
DD2OQp37JrLEh5HvkBbygsrYgJlc0TrsFUsEqR6bSjSdcdVqGT7u8ksr+Vd2WmB5
Oji9wlde6GC4WgyQD9rvW/1+GJlGmDBr70vCD7OiGI/UZh7nlt19uHBwSVCir6Ru
DiwWEa+HW4oa8TvHPeaRzBGqabm40buUdUIuza5oe5WXeYwC98GMgAYiEB2fitjE
OCqoE0okHel3tZ2dihWOxKPQAGHEOaZNPwCvNuV67onq3/yzDk3t6ulFx09lE+pe
51IlyXo9EUA+xSxTu1+sID/Oj9XDme0snLuEFC5MFDRHumxyz2grEVLVI2WugcR3
XrEzcybiT6AoLxPH3frNoQzoh/WBz5/n2nEyoaw7t5AJ0hK5GW8BqZH9TGebnWFR
DVjJ3mJAUZgjf7a3bs4jMsuqgAjuqhr7Z9Km+2gCpxORRpaFi7845K5WU4D8Wfs1
Nxzy1wiwWH5pgqpz6IJKJxd93FQQOYsVJ2JEIDpcDpG1zlxLmh4D5PrTKNLvk/+F
9zbk0iVjtgIP9qKQTSpYd6acWmQl/63Vjr75di6gvUmatpMLyWJ6aamfX5ikD0IG
72v5yyhtHoMDWcwhrwChkBG3yWvv65G+OIo1oMXX71ohSwuja3mqhK+meWygKPIU
j4v5RQaa7DUypxuuddiBOfF7mZr0FJLH9ocpq2bwOJlDs3d0NRrvqa3f7MBtUVki
Hxa3P2FIsvugAcN+CwyFUnreVuL29fLczegeOiJb8Ds/7jz3F5fLA0XmwzK9yYFx
2L52rUcAvzZEBwmvwRKCERp3wlvlFg99U4p9fCZ56RMh4mQH9jyjROqVLLX3pSO+
7t4hiXn8zzyRTKj/pFV1SAtaqqbnZI+I3oGogfu5YXNNkGpO+RDbNs1sgyFwZL9q
lZNXCKxZZ4Ues+uSN5yeuPhogM02yhonDUONJ/VDLHpgmEmDTEK9QvR9udhOPC3I
mCzs8L6RclObS52CrSoZ1nM87GGTXiG8H6wHr8e8fiKlvf67eFEZF71C+skF6jtX
e2+OvQKnwGQV1f9O/AEV3+rqbaSLhO67ELC0ZW3Idf5t0402i2VB8WoJ9EaeJ3qV
8bvGsTUyIl9oW+jqlsFM54fga6lE0uYw04lYoQecev3jn5IJGOtKjRNZCK2/JVeu
KKZ5/4hVh/QZd7jX1zV76IF14NOlA//dMqXTa/bhv4TN8D2lh1jC3d55o50vik95
LM1xH64wAkyoc+AdyZ0RiMNIVaCOYD/WDDLL82i1FKD6sFPbcKCYQYIDs/zF/v7K
ADW8WsUgDnEfwcIYdWfahUHxQWqvhwM8o07Fa5s6WQuJoiPztdAAOzZs6OSTbPpF
Hby5p7gbpwHe5NaCt6oQYbwI/LRAYqJL3UpgQflOCXZm3/ngPrSDU2C9/+O4WETJ
8mTq4gcnOnotxFwliyLCjAYaPr3auGA04iwnzfQacbWeBwBnGAtfQyDV1C/VB1d4
ORY16oEOtrN+u1vr8nCigmcqeRpSuLwzOaa/xccctRbOZbxU9uxcXplcPmvrJMeg
lA4QMQ0WesRzwtK3obLc32/W45JdgcfoEM8sFAvNynwRL4JuPYPAU6tBedHj1aec
OBbuvLGDbWv4uaZztPBmGRH2Hn/MOg8+wSVgvIAzugsRRTBMoqRCw5jamtHrCvdV
EAHhZYiSTbQhJZOCcR4cUmlZxgYvz3+HzrECQzU19rclRsmHAIdbibr1EBK6uEOj
lOP1NmS/cUkehZg2d2IzY+okPACchKPK4D9z2OHAGRcR1kd/cvcyhsYyfNZnTXsN
tGh79AIn8LwEMFsncPwIUVpaQYK1+RFnsysSOUVcZvrJB+epgMzkBbxowZQgfmiu
WFWpPEIfYoFhxiiK19jV/FjKXt9oJdRwUafxR6BOxtezZGsOUxmFKR8MT+wzcO78
oGFxoWwhNMn3kA9MjJCDqwcJ7L/Yen7Sq8PXc9/RGOSiQ6EQ+P4VeCENDT4z+1za
qfL0RmatHRNvvJcgRwAOyCQhjv2E5CSAgpRyiFFnZHtNEgcqf/7NZAhYmbeQMRDF
mkR7u84rHiDl2ug27M98jWOxRJ0myRvm7fvVtxKbmLFi3SHw6V91UpLd6SyUMEgM
Arv9DmpyDr/VML1iVpGbL788oe9EjRTlfvxYI6GgwMpgnYF1LPORLeI9vAD6F3bc
CGEWfGVO2aeSa34qsbgybj5FOJ1TICHHMywPBY23dmpAxUFV/4W1W3XiPkWsHWUo
M20Pf+NZtUGg+wxS1DEGjZmcsREuvJdHNtE6n8fPaJ/5agWtobJr3Zik+684bQrr
yrilj6+nkTw5aCSJsJTtwchhd1eFKttIgp1Ps3g8LE/BFE1QUAPH4SR/eQBbW+rh
bpRqzV0PgdzM3mnuRdyuqqUo0Tszv5m1Z4MqtR1SjvgJe+YxIGtaE1sJpt7h3UNN
mxgZO7KR839oYimF6gM0Cnefdmf3q3An8UTlZ6XaUDaA9q8swZndf0axBTHmUsaq
zDogcmokfY2a4SmQVwBiKWWnXEEGoBL/bcYckMcr2TzCeeUmJIfZcRSSX8uHQaVc
jARJwSLDmRkojVQ/Xco/OdXp60eDLweFbarHCCbM6OtSdrbDEBmsz4jAhrm9NLsZ
1i28v7YZ5WFXG8kKfJqvCobsWgxZIPwHta/3V2xco82J233bA2CSCNTRmTSxFCg0
I4obtpMDsHLf4tn6h7iB/Jw69EvAfK85IfJ3e8yGSvcOTfnXm9HdZ81qtQbw7INo
iB6NDnDQ5P5dRB3hZ9W9j+8E3Kwd3j6yU/mR5l+jEAeTu5I57z/c7qbUpWi1bwLv
oFkPudD14YgylpTKALsiiozo41CeDa/R4CoYkYP1MrWQzcpeRoFUIddxDeoA++g0
cJIVrLmVrAR3XA+1etgZS7FirzAYAWNj6Ya2EEQM0zlC3ESqf9YJW/d/WgqZ+cYq
E4RdGk2MVFzC2XtH/GGGWgJ+Ve21+vb89nRB8ZHSL9Efz9kEKBexiceUt9WKivQ6
8YAgqdfgzReybJASKsnN48B86VKAsvd2vnpXqXC6u3Rmco6f+ABdyQowCuK/3s91
mxjI2BGJVlZE13ORBl366WXtWASV/EdtgvDMOPfkT7QoBOV3+Vy0oKIQOA1xxk5x
QJ6JPZ4TgtWZl2k6+VYYRx2AVBy1N5kq2ZRK5Z/+Uycf+RarRLTZskGM2bZPCyVC
dFF98YNJ68hOpE0/ZhudGeLoJYcNpz7MvXwnR3c+XA1cI8ogngFrqIxrKu7dqvqt
mTzTsaK5gDoekMAsptAf3xGNK4vi3NtDke3P90l5WI7aGeoSYuN3KBJA/PTduqFM
kwu6/m5PDX4U5Rx5BiEuG0i23HhtlFQVZQevZhn9BkqZNPBu7I3kcQiEYRbzjY3M
MWiHRIM9PkdQz00V7P1TcfBCrBuk7D5fXxozNlAMqA8Cp07UJl49O4RG7RMo2KY3
+O0WOwag+RwfHjYdwCUW1ODnHTjr1uUdDpfEtTVo7WvtwEgiwYlwN8eO+X1IELUs
D3oshw0c50QGCm7L2dIXzgLINVWKUmyzZUFThzncWQjoFiL/j1PFWpz858MiJ71L
eSWBtrNgWq7K+DezDjMtIPNbDojlXZxlJyK/3b8TRRKIJjNKMEiVqFzgTChUb1Xy
HmQjzxdpoITGjxbm1ddCbIcpA54W7QC5mkU1EEXNPoZqpe84qKKqbgpnsP+ra42B
9abs6XRpmk/9t/OPQuByXJC/Eqw4iT2srrwDDUQJgrESwdyayNzNrt7J8H6EHMMM
hWjKMnwW7axpzQaj+O5AmDz6mJD9sA5FO40cB2Rxk/B+9nSgURBACVQ9/uMrwuL/
foARMKM3AWLwuOWX3rIwlIpfG5HtgHQtVU1Bsi9fr8q0br7wftrkKdXsT8ToLQSN
+hRtcpew9vw+EFfK+txUGLr1w5pRhVIMhwttvZ4oyfL4C+VjuxArmC7Mp73tbSlg
Zf5vKSkFet/FH4385PeLC0oasL7803C19EhyI6x9dE5xDOEYPXFNXykLCsg1D5F2
rL5S0TVzYJoVb3NhhqMNHMXAeyaLHZ+VJAOmDEhF0t0wjIccMBguCyvbUHHiukib
Qqezz7EnM4a0EjjqkZ53O7GAlRCWF3Q1WFFB6L/XZL6k1/wUDgN9lXHzx8hosN5F
aLzDgjdCN/RK7/oDguGcdtr9NT0RNPI0OCG0fnhqPTVSMgzIKoaaXZOOyVnxmG22
WhRENVkPaYp4nz2Wximli4emxeNaVW9qfDkLpX1sGDkcinM1spj0lGDsb280Tcmd
GNDKSEofKPln6CaPbC8OmK5EjUShUaWvNY3qo3aD1LeXBYn3nzHDtKN9aX5fDN5d
EeaJgUqo0MxPKUfw1yy6XszI2HGes+1eqZK6M/pQKaZ9iE9S0UvBm0p7MfTr2mW3
WiUez1sXlYw7BDn0Izk0z2ZCOQNm/SstCxzSGW36SxF+gzy5rflipXndRhKO2fgT
Q41caF+o/7DyUcdDEhlUlzymbOK2zdXbSiUI9XJ7p0ZyHCk0AP92OP9Rd494fbbc
0qGOdvrP6NUAT79iodQvPusQSzLNM2QFBOmHCtNW4uHz8TTIEt7Z9whCfkmyHs3y
m6wWyHNUV5hbwnRFVoB9foocEmPyxyZ5V6DqXG5P9fjgeqKVlD5Y63nssy/27uFS
32ccXS3AIIzuyfZAaMYDX8fmq/9igT3wExualby3hTzIV4IJ37fOk1Jo4GfBmYOW
yaslV3KOSEK2h/zWmwkU6If9qwYI4VnvhXOOhvOMbhMoaClAXodlRC5M7jdAd56d
1GDyuWtVqj3IInfYyEtUfyg62m3Z720XuPGl/3VunUbOM7hyaIwwSq2quU1Hq9qj
0aM7Fj+OlZnXGqr7Db8DH77VzWAeYb8zj/ZPm1U9nc1z0/NOcNavryGRI5B95rGx
ePY5tgbQzTEWxfkPAZjhUPWDhUDAqmL42ISLMd3VKREX01pJ/PBSbUJQsdqtl6Be
rRssXJgcFFgjSwQOv1hFBWv7dhN/Frn7R+0buJkJebA5RfSr8voQWZhDu4V9z49G
cHsm2PIDuzkoeG6Lh4/l+kS2FvL9o6CEuFA4O1VhvoE5J/yEbf1Qr61gCmjiJ1uj
Cxjzztva4ffhR2sc9wfjqIoB6f/NsIPpwt7fC951rqSAjigRm9Ot39jy70plw62A
l05NTdY7jabEk1OXOkQj9wbjD1UCgcYngXaVtpJTBqptIeIjXZx+tMHtq+G62k4X
1M0b1b8GCr3v8t11c6ZRY1TqPe2T8oCd0PX8hdRCuPUEKScOhljDLoLxEfic+5uO
VITDYhHCUYJfdN3vlGYa8cGe92TR7ObeNSKo5NUOgdls925xjxYPy4TptnIOrfqF
w34La7BHZbCQYFuRXYNFX6pzipe8BTZZjx/xXirBowvyVLYGSGilx4QIOr4c54q4
8UW08PGx/J8piv6+DjuaJwNHtziR1jZ2WAi86K+rl5CUCkZSLVtKU8p7Xce8NgkG
F4RJX/L6weREGY600suVHVMJYxzqoz/CXXkhGsFmXv70I5O+G2SqQhI+AX/nTo1F
gHgf9amFv7j6HFmEhY7JzOaiPWleNvY08SRXl1yEcWoH50ZrFdLY8JDDmgzgfzbi
3Y/OTGl7Rb7CtdGDVVW7TYgcRVZ/8sMxjT2RsCCxHJnrO9cjbhKeGxPdi/uDDT5A
wutflemrL7dQal2KOfUL6FW7iYeNYu9/ow+R9E3kvcnSN2pVOUPOhtwI6wOphNeM
uQ2nLTLwz1R2cxkKCKuJfih56wBeLEysiX0ixnOJQZfl23jSOZ8tf5Qt4veHsJBR
8z+TCxZVH88TMchEH4Yt3mbSWwck4kTQyVK22a3NDov8mNt/J0jyAA+MB0gFnn0j
FYKUOhQ8QA1gYU60Co/Z3Os8+FrQVQc2jH+UrwSo5hVq4AxO6mxORL2u/jSfFbpH
l+8+dZcetq2FBONnEGWOpyvQhovRLBD/TymMmFKawKel6a86F+ldZiXgjBuys7Ak
tA+TrYT2wq6pUHKgc54zxgQjbBbDrpjaNU0D+K7D81lrirNhimghMqQbZ9EqNXaA
2kjADODGjcrihjssTXW7irpJnPiOId0iBGPMVTl9Mk4au7mXN8o1z0tdygA4oMOu
W9ESZC2WdaH4C9SA86mKKUtxbjOI2bJ/0W1tLMoggjTmawaXQQ/Jhxgr2Sj0C2+P
tMh9Wy0vDfjz46ytQGILQWkdnmi0sfbvVRoGmBRAanZFDOSxTsQDZe5KFV9Exigi
vQxcL+MkqCNyAmJJvHIrbK3r5VxNx+Bhw9Llg/Fahm3ntYTvxhX6KxLtkyyD4E48
6FX1HIY2d7O89V/VjYKfQ75fGc4JECkNBDthOHZljHbg2HVJSMnloTcoPwx2D3SX
BuiIz2Snd1CDGBRJne33bWHbRSFuZN/BPbEKlA0zkmb5PiPv2zjz1L+XaTjHU6fE
Og/9r87DLcMxzv36fbj2pS7cLjQ/iNhwBt9pU/Y4PNbmOsAqqY2m2pBrbpl98aHU
xqvYoA7jTWfGYGrzMljtQk86q6zhU/q0S+t/Vk6H+HihdwoJm4x4lADyhvbynPry
XUseGhNWhddCwEpXZq3aMCaNJWh0CatKxNjVvA5djFl9crv3n57+Mk+YwIkPDrSd
FlK6NB9SRhbvgG8NWioCjclh/EtcIRJzr75qiXPkFy8c4Oj/nmkTd0Rd8s1r2mgy
rLV8/EpwZ2KoQxMDcklQGAiUenFxC7/qJFUg27tGUUUBjgYWwp+SSFqNZrM5SghG
gdJIeX11V5M+s2zZ3PsV4Kfxpn+7obwkSM0Na6WWjh4LiDXxcip6TUG8KZJ3OZD+
c77JF9m7yN4p3SWuzK/uVrEL0Tq2O75tN3FxUePjunHssFdCeM9B91VAp9kjSDSO
koVQ+PeToRAn6STj6HFo6YqMoT1aQqNJuNElDNBd8FaG774FFzZxTE/J4i0Xn620
zdVK7rXlsZw+YD5vzrtpTMw0RZxlASCCqgcfOctKKwSpfvCk3+/mqc44E7wYJSd4
yxZWVkuSP/NwpU6NnAn5SiM0mn1skATPh2nxOr8mh2vEloQWEjvsRGdPvZlzyh+w
3Nx+49e3POmmrRC2NP/S5UMEAtJ5YZkax889qYkA7OSMYsIZAsPVj7F2lCMl/B5s
IymBY+mtafuI9VgyeZ5w7lvPux9RE/u0iIltD/9R/GtIfw3ZUD84CmgxF7Aw5pvj
btOB0ZEpjRFyC3gIlqaooD5ncGLwnvzLA086YvZpPqEWwIGStmmfwUTSWdE5h6n+
p49UydpRXF8HO3xk/9JPbXJJP6r5RiyJNk1SUt+79tPbRqdDki/x+clElzheB/HH
YzvYXWQp1gIoMp6g07+HJG4gYcZX37eat5ombHfT9Rg1BsUUNtAueoUFKzQGEwu/
35aU0L1s8dY/tj/iJD/qO0aJRlZTDnvC4EFDV5ffcTIV4iyU7sj8kvZabEFJKBlJ
7ytJtD3inrYsh1cnbRvvVlFKGfpcNGNjarqPyU8UpKbgPOiud2dFIRSH27SyWyFv
gLaq1pCSsuwFXpRS7CYw6NAwjDEHnEWK0P8xZHvC2TPBfC+ChdYPxtJ8VMg+SvBm
DwxHY+htPlM0JOrEZniMHqyuZeQiAymJ+0YQY0iR7yLoHPpiX2i4/sy1w5GwgtPY
XYU8/5I/UiozrV814cGjbBFKfrbbDiBlsdZwYcKdRD+46JitGG+XZiCY5cii0lXr
HFXIkH8vBLC5ra8zd6lu+mydnwvw581IPTvLCKVObBbldt/EF+G/+qviZEBIf7pa
IGJFdibD8XIZroI7O0MWByW/MReykjbdsR4KkikZVwUOLQEW5mtUMiykQ1IW1xhd
j3J6qf1OLskNms8ZRFzIQBZMtOEitQFp0bCkctBR8zyMxRVP+SW+ZiBiRadYgiO9
L6Cxvr5QTs+R4aYeXQRHcsLGAM2CIm0EsZnXUl6fpc6alpCeLjBlB7ic8B9CFfKe
ZstVNRWAcWEP3ewGB/GldDN3dxmq9WxaI5SWjTm5qSLhi/zMU0RyEAqiD51yXdyc
v2INx8oJlZxdcC+0dtT1Z9oYhZYbtZEEkri7TVqvJ82e3jFE/HhL/0q2/6KBSacM
0VWgE9DZ+ZRRIDvt0wWkmuyAfija8E3e56M5wiVCGkKZOxPfZTo/HoElZ7XZLcXt
78Ui5vIC0fIRhuuXh2Wmm6naB1RkwWODlNK17zA/+Yk5PPRfVlrXSrjjkvykrPyH
2ABKl09bnmJCCmZVnPiosMT83Rd2rdJ12QPHMVb04k7nmrhHzcygnnO42L6pTYZj
xZ3t2IPD30KGuNxm2rfcjHZaTE1EwY/ZPgfwg9UNTBV0aQZlWjIax4xgA3aetqE0
HH9SLlA99+HZOLpxNn5YkYdkoE8Z22F0JKCFZeYmqnE1LS38uNh0Iw00Y2L3yzdO
Hna+GyRmXuKgdpO3vXqzHEOztj5ppeGWxRb5S6eHRbTElbQHZcoFdWqe4XZsnJls
Ct40UxF1NHOosH988T/XyL/3QZ2GeXhErlzs+Fujy8SPTukNs50V9HQOGoYTTslJ
y+fd9zRciY//PGeUnbJJtCMpcE7vxk81v5nfECskAGyU2RadsZRgBRT9c8KI5r6u
n1sEBjwYCh3CXmDF35Zjh6sHq48kaAzL45DCiyhvnXX2ewIvwzEwnhGgH4BNZJco
CNHekVkArNllqyGsYyCOZN9g9x0yBibRKZT3VB76PNZjsAuFctr0rXjPB5WCaS+y
J4hd7khHBdY6igEqfVtDtvsXVWGWgCfRsYW0vTFq567Iz/9q964ywTDp1gauFnns
EedaKXiG+0POnMqbMYPkPGNG0nIRX/EZHZPgQANWtjNyfFevAL9fCVWUO0XLBRjI
SSsjfdIOjjzTimiUbFtp7rzfTUXinHvLN8U/tw0/eQuXzPVoFXVit2fzMuz6D5a/
fK2qanmVUs9CyJ9XXNPVgoAl0sVyhQS7BkHeHcAYRsMCDaWw6fcmfoWIJPOeASBC
l3UKH1kE+8mOV8piR2yUQEo/UmiwgnGR4lXmgXfQTv6n5NBbL6er4/pj7OLVOM2/
usE+IGhNmL2/1ng+AOxiI5rGPxSZWBJR/kAQzh58dqDyEmsBFBfKPFx58NdMLOAq
63fVDCwYNsPIySi0QHzcZFUnB0L10q5KxVnaHgVjnPb4YwVksQUWuHynqmJJNceq
aRNVe9M6y0x0OvEuBPiXjM5B9piLPiSv/b9SrfBuP2papM3uiLdzPtwuplCUraT9
pqrarOf0E7a37SeXDW5m5fuUwFaRSyVCbIef3BdccO9qpMcX3e7PBEwq3g5qYiSs
TEb46qj4VvR+SWlbxdTwzwhoqT7W7S5Ufoy0gda1++Mz1wkMmIRUYo2gKImSGfEU
f+Ibm3LQWguCHySutkgRekSOxgS5uJljDbqiyVmLrNLINoM7pYeZ1FbtYzrZBtXS
osdEGSX0oB5GvDBfJOF+xI1KSLRPiM05vH59xf6WPJcyw+vGHOT+TBYPCAhBLobV
9BSVyee1tWUs9dkZYMg9ADeDhfLzfkNsftaABPLC4D6kVopkqDJ2O+FtegdWvuEc
M7GvsaVSjpa9Bop1A5XvTgM0VEZveMf7yuiq7B0jf4nwQZr45CcVvu6F+3TRuhzY
ir5a7cjyHZcI/kjr7+L3xzqzfIKD+qni97lRLzhw/bDfMiBL1SAhK0CH1KmWj8ey
mCPYoT0xMGmb3qud/E2NCnvpDKwfY/Vc6rJfeX6tH7ItAAB6z6OOA5BsxREMySHc
Gb2/a9tdxQEy8SP+mU3XptyGDWy01T3DCJiei4V5BGFW+YUbGeU9yJ5Z8Z/0RyxH
bJkWUTjeVrZ+4Ja7ogCvESQJOwbc6MRSZLK6w/4chUlr5x4cz0cAq6fMVblDtdXQ
G4GLCsGF7C3nj65jtCVYO9Nky49qsrE0r1e5obp+upgyCZusxxxjvDXJHTWCcKnE
St3vHd1Sz2EaVBspxRpqfYM8qEkz0muOaBFK90xmHJtGmVvB3ymmlHi22kJptVni
qM+9U5H4d5BC+jXd+8vuq4A/fCckM+Punq0XFmYcuZVnfLmP6T1HmGKXp9fGe8Fk
bd1YBMXaUehfp/zdAPw9JGJ9h3LgmKC0Z7JMdf7a7YrMzrj7FSuialVOVNcfBReD
XiqzDcSxtvkGT+nNf/jAe0bpm/Aw98JWv0iCie9kGZpnPOt0/SJk9wdb5ebfV1sL
nq9ulOGd5f0uXeQU1W/pmyugZiTj5IVGxFB/KThAFsj6d8Eopl0j5Mv/9/hJJtiI
8KMBjMm9TKhgNuf/ak74CWmv5cTWTcIxI9PKRQwuQ65QcWIxlN1De6AGnpLEekw8
VTe6MrKzbqw+KSBo2BYh7IvQZUhvmR8lrSlwlf2+37qrfIES9SzDBUZraYSM5dV3
jxQlkuCp2T60RvJQaeUibWy2dbu4yXgDjceogRz+/pyWYswl9Wcnj+16rKSgQCKu
w1ZPB9pglhVENOatTAjd0reTQ9v2NVakjjrk1ItzoJlXuJ9HP5B0qQJ8YYFMqLRu
SuJguIyxBvSNuEuTzw5Wxd3AFP+hxriHV2r09dof9jpntvx871FZPPOffhEsOjtQ
KteVgGhHRJQNQqRcy+3pv1uLHVQPoiCiyjuOOQ8IrOPXw3emJqjfGy6AYKCfumaX
RT04fZcj8pPxdJyrLc0n91/393SIsO22+dlAyIJ8o5/h7FPhTgyAbsOSBECTTDgr
98Pm2AiIh4u86QiNaRgcWcrZr9PSqmEOia5bnUyRXiwTLAHCs6ct50sewGDkbBEd
bP+xMHTB1N7T9MORkCe6aTYT3LmWUDssnPHHSW9HC9PiFAa6Merh5JWFt6tvTKfV
OztkC7yLRHjg4WY3WhNx+IP6AKMZ1hY6kxTFcY+O9XyGcPX7J3bKxt0rycoas53m
F12b08QnlrveFkZF7xBcqsoHiHV1HKkKL2grVZ9SRgYsWVJlz6kP5uUioCjBDSky
fEr+wyQywHkd1QMs8mqQ9TwlJZ2fN6pZxwrhUUfwtlqfuSWV/su8jnLAYztcC6b/
Mo2Z3igB5T6Iui+dFKE3ssLpaMYszk5U9akDxzhJppssLMLQ+t8zqLMycMSauKk+
EbBSTZBtbNLkSFf5rMZ6J+nSOBeYHKSpJoifGArOVStV+2TnBPuzY6sYaXayy7/W
j/qz7ZyqvtPmCHiP9o/CRi38/25if187HmJL6Z99l5LCYqyzqwOKRHuG3QOPhAXR
1XAtGw6CTWOuXo70M+Ouil5B8LJ8tjFgTFWt2+DU7w9ScQOSWyZFRaPkY9Ncp6o1
E3MIfkqH6ePc+8G0Fc6KHXzwBpK9+Y6ceQt9N8nDo3OnRe7TZp0xZaz8bFl6EbW8
EFpty7SifAM+UV3bUAdMUKJ+kOu6N9t+yy9uIWk3YgOF2I9Dn/3Q2GhzyPUi1xQy
ubr+h/aR6F9kIcUM7PPFhHEEdzoOEsma19hBmiACwuOJoSowgvaS8xWLtzenGEUq
mmJSxnzWOgXFKjSSG8EQCmwEufEjCDt+rUNSPNZS0DyE+3Ni1uLolTao7FBFRcYE
5Qj7xgAtFaocO6jBB2kKajVH9++dRNQwJBvJomnKVIs3w7cwFqff3lgTaQOgC9rk
WxbNZCzFlACweiF2VR3OIeNQcTYPRUwuGr67TFqRTdhJLXkmEoPnVKl/es9LuDXE
m7plPjy3V6Pb9SyDcPO1nf6YuMTQiJZeP4zchEj7UdgR3SQmbYV9uQSpsPqnqghA
0XlakK1TQktVquIE/iw2iRc8ClVNwwfFdoZb2Gyjr65rcUox/AisWCaZ+DbhbTkc
NJCsU6W85JxVpdVJ0xfMbwjbOluELFyQzlg8wX4f1SLgMejKRJjBnMaweEidSegO
yX7KDcls/oHxZYvjhxnjUJC16xA8MNWKp4gXeiFB4IeRLs0kBlxKo7cZF9wgiN1Z
IhsWJ9nD1DIYrgLjwy7q4D792ty1zVFheDVkG4YfJCxRcBBsGa4zuME8qe1BV3bR
4bLST+rhy1HNqWBg7ya4QAU5ZKSQ8+mLXUhJzGtHOrjvQsjvVttX5DxEQsfKt+tQ
cfwXF1qsKx3UJmmmiX+GUtDbPbyr4h7qslsHZzC7lt2ycJxDjyeN24fOpFgwJnfH
wOpxb6PesptTnr9wauR667V9bERrf7KYuQSxwOJg7EwoBMPHwT4ZzuqGOTEve0HJ
89Wjj63t9sbrJHhrV9j90IVgbt8UIYuJwjYveo2j/wRZh10B/l6WJqlfTNOb6WTm
UGZuRfKOa7VHZzTZaTH7ROxGPvOP4cn2yT0fzkR7x460s08zIR9m5imx9ovT1ALj
AvwD5xQx64ZxqUBaX1HQ90ULO+jk/ilfV++9LyTOOpoDX7FUOsRd8AjpN9na0YUD
MKvNHLARXHQ7Pd9NWeTHIT3Auf759hcL2Z8DjAm7hRsLajLiXJDYCUZB5l21zr40
6W0vmYKnq7V5jbRAvkozzYD3lbzlAcYYjWMpaPxgMQkcTmO1ulL5vmt1BsA5F2nM
ZHezIk9YeOFNhQtcjvy1vjLifpPrKAUK9knqSqoqkuKzN+/3V1w7vgMJQM5ecfHi
M2OIrxhoRSHEONuUphsN/460yJp2DWdJFNQRas41Hpz96z8vwWY1fhR8IQ/bAgKu
bUKNFmwHBag71nSYf9Zl42FP+fhb72pWGDoyqG7aMrMqWblpcYCfLF7Ua7a13f6G
A6LbBB8zOw/qv2OGzGcWmw/uTBmHUkW8xOgY/hQds48l1DvZ6U+ruVe+yYD+pTb8
Ml05InROrOnjL6xNogCLfFz6xQ1Boc0myzH4T+1UUC2X0RqdVHzIJ1/U8ptPDgLQ
SfATNdTwDf1GCCJSSPNGC3xzrBNr0vx7RjGW3I5bv2opfIkBEH5PjJ6X2O5HA11Q
DC4KbU/c8tlHn9BgXXVXog91Zt4/40duw5Z+dSvlZVZ5twheuLlTM7fbwou4MAzn
haUgaFHrRjOiEBH5OAQZOzq6ZUK0IeDpzfCpGVnOMo3J6Dp3zPx8O4n9M8ja/YTQ
xCHFVMpmcFtRWaWORhL6pYgSZerlQ7VBESFwMbCKOHdK+gshJrmr8tX+jBpHkpBI
nhRnI2qZIF9D1BkXQVaFpMJwdVZ/tFa1SmKPBSVGLQb9yxH4TdTlTDQh8nCtIlVF
VrIM09FiVTpmBPfWTDPz0io/scwSBhD1446e22NWY2Liy01+ky8BAddu32ZF6dbX
VEEyd3B4ik/WhhAK6HVbc8TMYAVEeTQGjkn3WKR+fBeH8Z5hrS0pj6hWKuw7aC/u
HdgWIWFO8dEA8UjDeLldrw++y9+ADGLuQlrzOaEVRH+qjj9l7s+rVKFX5Fn4GLDC
+6YhVVgQkAPWQC1JcdkYCYnw4AS8DsrUGHMT6DOS8u1wmTuSv9pBydYCFe+0ZAj+
M7kUiRVjRTV96K4RgoC5DqpNjdMg9IlXz5b8gPqWvTI0vkJfRsodLx9mCOWdoumY
tvP0Dr299swQE7THpfD469o8f7BEXSfXA8116fHk12jfPDV9OeoYJINwzGopgKC3
qVv2brdJdGc5hJ1Pkiz4zlbMUD6vXXmBU6Jc+He/TXECLeMq3apbD7B/kpoz7WCg
2gFYdmbthUC+tECyjzKXhx/OE10S40C304/9oSek2ShIhf8iZSU0MJ1HOzc0PUyW
ZeY05Wy8RlwqEocHiO3FSwFQCDP4SMWwMm0FdO4c/oHgz3yiDSiHV8/zdTOpbFaZ
PGJ19SVxKcxan4xM8lLhE5D9S3nl4TEnhRJHIM/L/Ti7JRYI8dvksE4uEghX8iGN
PRhtzynO9CYyNWft5sun1Q1xRTffBYtJclwXD4MXdtl8A11heaWx4sg/wuYa7S2M
cMnJd0WB7/cc8r2AY1+PNyTKzKuBK+X6sL9XErFkUjTMsuDydv7H+xc8UjZlGhI5
/hUua4eqZVb/E1qsZJJIg+UUHorjwZNeh27Ir1NpVnoZvyIcq+psBbTdRLN3qlpm
cCFMiAqQtsxIcbYbiqQbOJIYIHzALiDdCbwWx22jHQ0RyZN8+b4q7eJxRa3y+Ia9
R2FYASXRJNa4NeeXXL/B22dET/+tRNBXh01bsqP/fEbejwQY9zlnkz6ql4zpkxij
ua+HOY2j6SIKoPGaJTzfdmR2s+awsbQmu/Z6/yzJ7ObJhpAXJxvWYBcwhql9x5oB
edp7I/DUq7JmvxEBI1Qi73QcQXAcmbS3qEopGKuVp3o7a3ysKsktMp/18UnVuPIY
2Dpetwr1/5jAIdEZvqpPqGqXG8VIPSg1iQLVL4OkIUfTUTJsNYJWW19dRP3iHcLT
EHBdX28PbbNL+dUE2vKA5KKY6icVPSFlSb6h79NETarz9C7igDEw1EEnSELtWxul
8NQtymjgAh7eOs2dZuzHQtWa+1pcCuG7KKAtDZbsJfW8wdW7ZMALSHPgJyliNLLU
CQUi4ZzWl067d5rtttZruIOjARnOLS/3M/pNewPP2l57b82BgsDnlNm5mlLLGRb/
OtSHpRZNsLac9jT0nUtFQ69TqsoIqowsws9rKlO7GjpRitKB8pnmWO3YRjSTYawc
YhUvTp8PX3O8GW6VffxAgdfISI6SYjJd9arfWauGQrcBS5939Bw9QMu8B71buYlf
VttTjcEoddxnXzTRcgS4p8qCvivwJ+u0gsWWigzXb9NllN1AJ91x4Aak2Vfmg03i
AIFvwbF9ggqHWTyCS3Z7cy2DFwDFfmiXPYhPzx8aGy4P2OklVHkNLc/PcyzkTlRk
p6uZi1TzWyOC9RysK2kHhkZLnZ8tUXZA23UiO2BJIqACEFgpwnb+TvYhRRnsTd+V
hmPTs4xEqmbnuyTcZ0Y9OMDD1smH5nF8/Uc3+9lXAf/8kN74lyxwaX3c/5G4XYYa
779tX24y3kLHmAYwBxPG9N/QWlc04N0tTPuWiC9TcH7V6EHT7+h9aIAjLxZHB28t
40kXdTbc50utQW5YHUrP8sHij2ipuiO4sNGFHyTFEpiSg85bHUQkHPvB4dqqDOUb
j3yKHKRrbxp4Ju+K2XyboYQLQ3solLY9DxYca6CVV3BStv9NirLFqhRSvLSTqO5y
DxlRJeiapfc3LkyFGhd6HZncMYiJsnMSJSYQEs/p7oJFKQ9m6T9hTREcN+N23OK5
rpAObJRKxRbH8g2ltWYaAgN2nnqwKfFgoH+z7vmDmwfc2AJjCk2o1bQKb8OqBarq
bPFm0fxZbU79PRhURgORySFihuHByleRfL6PbJHGoL87cjLQdRMZhTzqK4/2N8qg
JLt9ZKsrzs0eeQSYsbPknKUoE2TspTaL4uTxaOVBFfMn7MEbDbbFSMYZYJNwn8DI
Rh+JTA8050r3HK1siSo/inl6HRsL24j9WTwhC9D246eJOsxDHKtj0+0Q17OtUl4A
WPuuxP+NNyh3qA856RfGPKv0d1tzE1L4nfGeB3+4aBF7ChuHybxFiXoYlHjMW26u
uuupCm0qdJoEu4W6Gl4pD4NBGraFKbHie/kc2x2Bkl0lkkymmgnLnrbsfGOdj9CS
xFq0nw3gPt9lsfb0Xtje3u0mU8cslHPPeQ/iNFvqOmBRlXxM4fbqd0A4h1tI9aqg
LU3GKyNEjKA5nmmXd4wUnbgB1Tq9bGHj38P8KA+Sy6TMz0ohUmBolXgbLMH/9CXP
BFlV40VIkjmAA4+z6zB0ZDMuHi+2jWf2vKITu55dIAGGNvA2jCv7Vxub6i3akqkZ
wyWTxWr5GhGsYHoSoWHgWmDdJzue3hJygUgr5rRahk4NXWSw840fazmZBY/aduoH
0TAZip1NzPCZJWnVKPj+EJuVJGVGwOKl5bpRMpuBNx3Px5IP6jY4H4hWAgXunuf7
CqKzreujinlYze4vm1Uw0adjO4r4uGHQkJwt/G6fLkQuuripZ7U93cYYXHUqoa2y
qwZdT2LYOdPxmYgITaJ1ryG9nPpUWM5E1HplRi6Jv7d3XLeN4sxp48WzRNehfL4U
GClKD/Xdr0al25q+J4f2XgaDXroUYpm2nUifnpsB4zWANUhNnrY2FvafhgP4qb+h
CJv/y66U7ITYioNn//jEgGp4GRAU1kuEC8VIWY+UqyCqsAwd6wyu5JMLWXJ4dYt+
vj/CloeR2LugTap84fekXGQd9/lE6U5pz+NWjL9jQiVHZBewC15kPqMc7qn/E0o8
sgfRAQ6nTmhoVagf1sfzZfWoJeJyw+ZlGt7zN1iZyxKP9ksRp8y0mZxQrSSgXdsX
6EuUJP2ypdCxcy2pi/oziVAlTcjfqXR9AxyTPkH6tuenlWWF3xqJFDmKTM6X5KbI
PDtVb1MmYjr2cRJy0k2br9CP2BGZfMkuQZi++BPNl1vH8VDh4yGfV8oVCqhlvzTF
KZWdSTznPp2ubeZvSDs7m1jPNiF4XkewTiBd0x3L/IpHcKSqdQDanuXGzxUprEtI
9FMHxT1CXPcU5Ueap93c2Ii+xD+rB0KI2idUFRRhmnoF0mWiJ0QTMzTXnPi5Kjnz
WHYFisf7MhBiLglw3e/z0dtwpTWxaZIOgfBKbq4yV3BKGq/lk7VSHLm0VPhed4tu
aIhFFS19w8+UK6h/I4eTfCquuqbRyjFdq10dA8uQ4RoFOtIyZA5fBOQdYDOYEw4d
hh40HNNpYIwZCulZ6dYJF14FXDz6RErPp5qtiTmPB/yU0nKmZXxiE6GP7Ozso7si
ZSuL3nOowuF/kyalnpUxOWDkUYLylrkogO1Tfa07MEh4elcj3IYvXb4kL5Serf4O
9Zny+6HI6Dk42KLGbJH+ylcyK92Wc2/3hC+m6PptZcDoiRjGyAVU89N9YODvQl0w
4RPHp+BFffVytI84Sn7pL+RmLN6bkThA7sytzL6tPYnr/FviQuW2wxh+H6jpGxck
fpRTM2awF0ZFjjn0xSa3FO0olgDocdLCZ9Y71u7bNoHN2WCmIE2ELrc00CB0nQ+Z
GX2MkIBdB/Tyayvj7OLjLICJ7hTRyXlwk4Hcno3pMaUnW7JRvg0z04svwyGIGizB
ZW+pEj6Ov1v8Y77Htd9jxOFBBG3qthbqfayNH11+lp+n7TVd7ns/lkyU1pGk+tO2
0zQRZdzzfX6UDdFHwmb0wJxVyzehuvQhbTzhQjG2WOsP9GSeYVhCGPT86JQbmyl5
RG7YRNMvOgPB1irF8WRXwePHJxMDrvxtnbQASyZI9l/QrcJem73fosH/cgDx2XBd
JoMrlkciRM7aksdwFb4/Yk1AAG+Svi3vYYCO46hLzH++Ptqd+c0fFgL/8PZqc/vq
DcLBfQlvgo2jCK0OIoP3Ohic1GNPNN/IKBiOP3bCHWrm+E2a8fiq4Hkv9zIXuaAk
LBfZUS2AxiverJBNz0XpfkUzYM3USqgOitwS4dUp8hzRXlUQl9Y1dxJ4DDmPYDnY
R9KUN4CeFlJX99shKPf/O0j/oUgp1Xc1N+kPVnr6sOI8WelJTFS8TscOM4U9cdn2
eZGicCmS6TeYZSw0Kx1sFyWHesFDY0W9i5ReOn7T1TIAEzxeL0oYEcrMC7fXKML5
Fpa6AEzsmIGi/PR1uB9K+4+pw0U35L23hV9UIjEVuJJDnI7+DSEpPAxGTJtEKz5v
/G+Ss53xvEEBoGuroNgbZ+xp1YqmRI70q47se1w3iTRU7MtlXyv+lLRS2z9sMguu
CsPFpmmX8wouy/rQt5tKhK5tZ4uVckwNPRavLD+g6hQ0J0XhM/skacePh7xQOZqq
CG6WTPM9H4bbR/vwDrX1+ClMtW+OfOOpONZtns84N8SeR+OFJfkuQI+0CFFFQMQc
BKwdi0wLEk6nKou4pzXBcTlGNsk44dYN++SnemRibN2mZ0Q/BH3fNzq/q75NZGZ7
U4hKNC99+xlv8mwiWThRwALwGuJ/U44n4nlJyqt11GXGwgdsGnAK9mfq79IkWv/j
IjR+CmLdDURRlivOcO7PCiM7tI784Kh/EITqLGqp7fX+z1+IZA4eaLz7sLpmGdz1
1zddiK3iqH55HUxXw3rG1VZIgaN5OTUu8w1bY4MWXiX1LLZ0w4jbjpuCAQdXN/i1
EyIG2bMXs9qJgHA7B9pVvljVb5Y7aeMZDkIneyr289Jba1vE6VNB+grFQyD/d0FP
OdQGVFUoBKWS23jYjG6rVougLjlE2u167JLUJA2eCZizuF7hwL8y5c1PKg+CeqrT
c940k7gp0hAQ4r+yd+UWe6Z3ilMOJJ12HMF7FYXZlQc2b6mRrxhGC2TyPMoDhCxY
eU1TmfMNshaoXw/k1PPHEkK2iKqX+o6BmsPFFRFLdbpUYHqDb98mGn5YEHylsqvD
yNFp0ycqqHMdJ6mB6RZythxVMW9UHJxs8fpMpTPXXZoc/oP7zW/Z0wc5kd+fkF9U
trwiFGzTc5H1+AjWxu+grjVq2VzP9LcnUd/n6Ge02/ug1+PaXMuNQpFYWpKLZZXE
dXdtG1om7mQcxJyMbQGCg4tJNZtrDvqGIT4Z5Xm2rDpnZwqKflLWu47VGU17o5/G
G77A6UPqFi2A2Vnw/YXQvnsN/5QiP+qOhRU2VFNz3CGT+iFlMjqjjnxO07oL5k+4
Gv3WSsi2uS+TE+0bcDU1Uy0+JxO5vebK0KSQ23k4FwBIP80paMqr1HSqB2BTwfVD
cZL+hkjr6WYxVr0njWFPkwkw9lPkZrZKgaxU+ahPkqo7kxPq4VMtGt1lmLX25ut9
R0uPwvplgFeD7BTnqywdWYIVI2B/gAlYAxUqIYlURW6RChY1P41XdCg1OkSvqmOf
8A402mF7hO1FmN/EyvxMv5/7IhfxBmmBg9+Jmnb2WUG0NZGTmwZCALXD7OxYIKAO
CtA8mQIgBgG8A2gFfh8XrJ28BMEjIkETeUP/2OTumj3ipath6hFm/oua9D7btm7w
hgBK24t8sJDIGdEhiMOBZ9e93yolLvjYoi0Tq0dDunHc9R4yLzsx8Kth+By5rV3v
a9p3nNCtBPVSGihmiLaubNZDUoBLqUogtCykvyCVnumNi8goKZUPxm7ksvUDg6PJ
fdz97B0XdOlNcUsNHXzcdJuo+z1ZF7/n9HvHn8DDMz3BRFT+oxFk5+HyDZ/Ybj8B
cF5aCK3DKOKAPk9wO8GmPLrH842/Cf+pfm8JW0nQuUOG6B0r94WRc9DlL3m1Aejm
ox+qPndPT5M50SC0z1VPw+wQy7f0hluTmjeKJWazfjREDdDu1aCpQXO0IKSqJPKp
CJPjB/xPPJCNQUR0n9tPRGRrt7cJYQBUNtgXZDpyxDaGMk2N8eRxS1+PS0gmnbac
yi4kXCoeRjC5ulNy/Pk8jkYq/s0KOCwrbk0HMxqVuXjFA3OqUdXRARg2dQkx7v61
Xw5TsR7Ky1PZmX1RMT/+WFYwZDMpkotGq8LUQ3nO2EKmbDhTD6tcF0bebc7Lhbum
QY3aMUJMdDlmdzBLh1OjBD60gXq1Cj+PT7nx4vqBka3YNAP/VSNne/x+HH9ZqiGK
bQG5oBvZAR5+16jvOh6ReicCXmtZa33tmqU9ea+Nxt048k8/fYcqrLF2IGMS1N4V
lEeNZlY7kY8PlLTHkZBvWFGmc8p4NdbA/+br5+gCAXsL+KB2AEBng3Ofy4ezPHC8
WKcRBOToYy/WvXkJbt+Exk19e1Fb7OjgsKIZEAyKoUdBj6Aa+G3F/eDDWqu5KwN4
FkODEXbVQJKYLoXl5bNnhQyVA1cm+h1IjdAIPZKCDkpNitONzMiXfu7F9uvujWAX
xIs/kCobKEJh0p1Zc6AIt3dFujnB22mIN/uy+fggVuzDtVmDwsZQAxJ4WUIH879t
ckULYmarb1zohtW504V/J4Td1FTzvzLffxQle/22nsRZ/duIf5OSoAb3PJPjIfI9
sRWDu5CP6DzEkuV87ADI47djt6waODdnxr0RcqJGru7GMavFCJHvyO8uf4Yb3upG
ZeZxPiAB2VTTDtPYx/3WG5qGh65LNK9VZIlmJYgSuCKBWR1QsU5czKZmUgMGmUTO
mbCEp4VKzCLwYlGr7nGfZabiwY0DJhxEquMtEQwwjm3NDqp067ntwJulzfjyDWiZ
ncYbSdBHWglBsXZ/Ng4FBAUWc79MlbvyA6n5TmWjzm2QBkOdO00JueORZEnYm37G
e1vjkzrdBQfKOwoMhb0sFsUwxtUAMjfWvA+vpQTAzeSN0SNDpK0cNn2Htcdt5OTA
f8IKeWlT5OY7vPUfSoem46U6D2tdFBGQRId25+K1shBjK0FdikUKl47cKB/noKC1
mItimfHxTV78FWLYHjWhWKoerTusGuGHZpLQSPD9Q/ssggNpqw088x6FmVZ2ufIl
sfnFn8X76Yw3lUkra/ITEcsHoq45Grx/cRi7l9HAPElBF/1Bo6g09oduLR72EBng
/HLGl0Ac2LNqNRfKweBzsglJnXf5ptlnmREpjKrAJtXC4FCR0oUq3mpargsgFFHK
wygKWIiPBFJIp4lexRiZXqpOJymRthRsi9NuadiazTLHkWvOyN5daolwqZJO8NBA
C2TrLBDMK9AYU+FtcEGf0TzhgoqAjEeclBYKBsoR3r43MGSTfWAfUv1nNQcbDnYZ
v59Nure3vRqhjfWOUsT2yqcpdELNhwtyZzwqFrXU9SCOs+bfLGtqo3VYvqLb0WUG
E8rTZ/NRQabNwB+eBkxStdKT4Nuh+jVUD2V9priyFNk3msiZ8vZ2XSnpUtah1AP5
i1uNAEpr0uHdDb5cQYocCji3jZKtvZvowvnKNhVuNK6tLsrBquYD8ocoKRE7Dfxp
uw9qdyh6E9rRJfdvTA0jpqGGIZrqGDRFXkQwoG9n2NpTSloyJjdkLR4dioxWe1dT
ivw+bpf+Es88NeZlvHWN/Bgub2BbBXHoRmrh8Ust+9WmYLsH9SkRaE3MiOWXl5zo
0EKyZwov466M48TCpPZw0I2SxfOoMkruE77vSuu8gRlyJrK+H5i9O301MD9iH22a
uhsvRT/kJ/id9sbzAIGJhjXWmgLEXy1SL0LdCZ1uS4Tj3AMa5fP1CJF6ZI/NCqSU
s25RswcXdkJ30l2kf2GrbGZCh41uz97HblPGy+wlirkSvFDjR6WLjdgkFPVj1jLi
pmkNz/vqoIkST/8/2rzDV9WOJrf8hiUotutFcvxVNACwGEoYXOfIbKhluLAjf+VX
l1uki3oJw/59AWtBdGLADom8eZ9auABD3oIrfo4flsiZViL4TN1EuqaHHHhcPTVJ
MxtArk/fNzavQc9yxOz/fZvWIO4SnndDQTw4cFXr2SyOzj9qpPFJ9JpMUdSFKEHn
Yhb1uJeVUwCijy9hENEBlK+T83YsSXwGSiefCrUUvNzcZ8IHIs473mIbGYtyeFPW
EzNZB63D6Xh8I951xEaiuH3FUVJssz9qPRHM8THSXTlF2bfjmyedSu93+2WPMa2c
ZWrSB6fGILve0x0ZNkYdksC8Wg6F6QYMZaXoDqJroBiupI+Caa5v7dRsxrJq6C58
BVoLCfNCYPPlBl0Iobpg9u2EIoJjBYPKptpDEXK1WdQjswiNAs/o1iKvLtBy0dba
D6/esJ4q8m3GHQXRRB99OODH5YVc7/NlDMSUlq3zbqW2XdSpr1hY8tBK8bF9KB/5
vvkInB4CPLVLSHtNc8eLl3eDzcLQ66Lf6xjKInflipfFp2UqsDEBSi3IUC2JMFgi
n43e9QVAMsNQMGDPhBMnbRuuK2JPtbGid8ZbzCjDfSjG73KnOQdvBWxnKio1CuZ9
J4OfBes4ocOy+//v0DEkEAPEyiwq7B7fTYvhebH92gyUm45rB3PVFB2g9pQqG8+m
26wffHcbYYKZRhQJWPuVMWhGkpTe6auezu/EFSFEnVGuk26cFa/h2SHcLxgF3Jfj
Av8acA6CkehsIHHpGoXMtw0d5m/T2YFDJWjSvfqvHlBMPEGidK7164GDMkJ+E45d
rbQ5sLgtPnMY1uwTm3XzWQELLJfGttjqNzgPIQh+w/qaDpEbaZTeT+ZBxmjMaE+2
W7uDvxaeUiaMr9PDrRDpEw4eHzLkCPGnm2fBVps27QwP4XajoDbLHfVDbyqwIpSd
gr8NLaXojUmH15PnX55YMwu7Z7d75/07bd3vINVL0+VZZ05P9et2qQv3PAi7KRkX
8+VRH7NqxDdjSTjhZZ8FfPvEYsIkSTPyaUqWr/t/uDk9bYAkAEbdpSRxyIcRejgZ
9bxSxWf5VrodSbND1cQ6IoFZLLOeXkjZLxoaPkGEXvuBka2gAYVB+HjG8BOdVIaG
3IN9ZLIQ+2KJk62nYMZnRL6+vrPOHCH3b5n3cp9X1KQSviibhKML0/GogGEdEwi7
QnyHZmIdS9mSpzSM15/pJJQknnVB/8p3Fzs4/EqMgQQ/erfwLqBPrJWDXwtFN6mx
fJFD9E0xALoqiv9LMo9B0GgoywcGTbCRqzUpRNWwOLO+kSLGGM7TreDFEfmqte8q
znWo8yn+3b9RQMnp1LVDhhz9mUYeo8bj1kufRvL5NvgDyTyaSuwZu4L43zq614y8
4sj7LbuoAacTjAaqz30vz+uTPbkzkgoRpalw9ESZ8XuUtuvTAOkfFRYCDHuugyVo
QiDso2vfLz7p6P4L4FGznQ0Ziuvlk3NU23GiVDytaqy86guSYP++b2EC9VuTf48G
WVerE4Px2uc7s6Of2wF+dbi8ssTlgIEL94KLf85VObtOhSiJT+C9C6J49+z9I6eF
GGsU2hFyHAmbrygQKeLFxzt2HuqObDtFalpEHrB6tUUZd61P2xlYrGZcNqyeW7Vq
BhiAl7s966+rAmVsENhEySAg0XFBa6u/vDhD27wKZYXeWtqPwrkQEsZgoN4RwTIc
CFkiaPG2oy884lfzTzDCpGb+K3TJpUElDsO26MqyoVlchF6ke26+DT0CgWGpgshE
aSO6ffkNVBOCu6I9zZIXG43DcrV3oogFGI7cOQ3LYBnyvWaVW1nokaQ3hUdj/4xM
ALHPjr5gSjqo2Q2iPTqe4NaRczu/jK1lBJXntnB2lzfM4elyDGgwm//rEj5Iajb2
URCAcqgvowHrfRnHqtK9ZHwaufpvc/IWHkOyitgBevVzb39/CEP5aaRA8ezJx5xs
zXeOKj3ABVSMzkYEpRUX+uvrGGufeieZC/r+eA15rDgebmr66sJFt2tRtje6ohd3
w/DDt6Epazk7behDuI+g9elPFWko8XlxjUmzV5kMbDaa3QACJDRdAp35S4dZgMF6
Lutx9xTobh4gf44R2plwNGy/oyf6059i4m8kvV5Nku6CGq5PO1W6ATjM2uL/FSxq
SYljiN34fO1sAKirNj7nViVsg4ICuXUbtGTPRSo07kFnceRAmZfWFNt4ocRaFrTl
W4+kSXeYk1cfNbiikBtmuslQ1+gzP3ucCdq9rlCRBkkSf76Kb71DOzzBqOfGqXRr
6PFglovT5bgL411jGtXyEdjpZLZLiFB18PdwvZzANVD5eZHWPeqdZfBRJ04bUjnt
ys5qjZtzhOzhlwEvKqIJ2oly0zTB0IBycVxsR5+BkI77WImngnvp/K2yH/pIL8q0
BcH9+c1CU3+QzKM0G+Pijk36T8TEqt+HvxqX9ptjjTmhx0I/pM0vBLnJec3kJxpz
3nZDMEYAww3vLMqzt0ODV1lEPudNzd4SD1QM92dGoX6Kq2u6eQa6If1z4I6yGdPr
2F0oSGTwr6vSmlw8N4+SsJnWcQL1WoPYnAi6dOwu03jYMgdgWPjTYvQEoph7ucGP
2Sa2oo3qSOO6J4h4twxkKa/vPhWbaYycD2oSSTiW1iFT0+WZsBdClQMm7+ccKo8V
DtG8JPbQVCymSsBSM5SJA8i7RpUG3HYtr27jLyjhUfE1g8Ymy7DQeScO1gMoawaP
r1Piq5sUFOVi3hGjIboULQLufyYuFLqR7wBbqR5riLD0pRhrBSrXGKI3bKruYTDZ
EbEZe2j88hcS13gl0s0Ayoi3wm6II7jPug0uIKoL8t51fsUVqyEtbHN0oN0IjsHD
DBN1T0jxXqsdqs0BVxsmRXRf11JmULyhYikYFAq8h/h+keC0xOZG9jDyDidvvnSo
2Tv37MHv9vjBCHz2MCIx7/hLBge3EWaFrGv9a6Ovd8Z4dDtJPb8Pcmt+dMT0sxTa
tsreQJwNJ7/8RO2AuJa5VoW+48CCLBjWzQ/ayLiYeV6LQcK466DZh4eIGWC0I3lx
Y0vW5+M6706Vd8BWNRu4Zq3aBE5F7hKPtUICUeYOQACXBBq+hFNBREEm/uyrA/83
A0W3ZoUWBiJMKdTx9y8xud/+vK4AN5RFhF9cFMhGN+mrY39zJLlbhDc3YycnXoZd
AFpdLQ22pvkyD4ta3YYG2Z6jnEjcy02PTEJHGgcRkNlmpXE53Dl281eXXjeABtYS
Q1Kjg00yEl73MAlGXw1m1/ijsbGtbZgVgSkTUqm7nt5iHDHzdf1A9ng94Oa4PlE3
fYs8AU9Z/GDoMoZSfEsB9HhRQOs1ltbnfsMTReNnFpHllQuQPuPVj3BXD9/rOHHR
vBytQnHPTBC+tAkLcYCeo/PJdbvmo7YUnh4MkpScrTtFRXWU+chOsEqjZPIU/7mp
MkEDWnHMdRZU0WRLKcr4+SFgsbCftbVXfQW2AJ4wb1JKJj04Kg2M4o+7D2L+E29S
xtePDLka7TKsPQbeOr5AqZTf3S3BnQ8Nx0v/UWiRqy6yooTZgsi5xOlf2VOgUCUm
NXF5gQCzRxlS4WEr4lWxVfLGuFe2iwZP/nXi6voBv45kb+EHp2OJfKmxJnjgfF+p
01m3lzJ9N/Xhz2HTNXbTy+I7Yg414oJH+EXJHy7XKJXY0/+l24tvIo2GhEd+4hQ7
Sx0nbWhmfs59r7/pglA+KLb05BfL3pT0NgKpjkCzWmg+InVpllubcnbb3CXicEaL
2fLvUUxKaZwRXKUPYDb3wZ4yfuIU2U4/lvxEnYDRqyBid/sn3JOvmttQtNeG8xwy
aSKSlDkpnSJYSxLjg2nHRPGd0opcloiyHq85bhUWtLkdNbPgnof1x4RWP/QHHKxQ
TkIsQUDa26z/hrQEqryPHhYD5U0uayeNpR0O0d3xKPncgFj+c13WTgWZKnbodYxi
HeEj5AC+rrL2Se4RsQVwQrgyhpySwAfawFTGTJwN66uV3z/dJHHWrBsIhNtB+OVp
Gepy6ivIGuWfaIwi2rjZYNFIATdmw+RP4B2FaleKNJ8iVxBn0VaLu00/XNrMDKtx
Eip+r91bFoUHx9vzZG4wpeNtsMpvECMsKmT7N6S/BgRF8+QdTimoDAa0U5UrOFRk
58Lu0RcnBEHpt+ac7ICp4Tr+9C3WjcGNh9a8q5A0dZ7AawgCpl2P8sFX5pAvZLz4
sQDz49qdg5cz6/JuhQ3KzTBPrRNFqagLg8ENph99jInuF/HJPzoHGniRIHyEnW0p
cCNNR+nbZr3TGvR4oDpM5U3X5j263EezYQ+h9Cqb61qTmbRNLkFblzNuwbOb5lZ4
jI0tzp4dGypJWqZPpliYs3QwfXr9UPy7VvqcnOfTNLH0CaIWcK13pYXuV82+r4MB
amSf+2szZNy5JRd4fRsWEdqPc++IXJWjC8gQSCJFg831s96fu6MX5CctH1dZ81Jc
0fswVMFRtehWpLJ2rnIt7VJSKKr5vbTcvyURb5hGSlNRuBxEpFSwJ15xcG8O+1DP
I57ygbB2YnLPefws7jipcyxJyJuAhPFER/YRlK/otn+5tLOVwsnUR5506pwHzNJu
eUoMeME0JgUsn+n9owYdiBV77VDOvw7dPvXivIAzK4mioZx9GR2xJsapDJiLWfK2
xpdMHvzjvJZMIkjpue3G74aYSKe6ZmpwBkn2/FRFc7nzKV8yk+5wY2oYlfX4pF/d
SI+HQdOqmVEIduqCx+TfHlrx078p83XM7DpZiHPjt986OVoLm4xM0kpDuLU/JUkh
+2WR5NfwKszhYlBjXjea2BOEf4tWbZ04Y8Zl8/GHdC3XjKPyfgoXrDErMJtrT9Ho
sKyYIPFKdVDg7KAuFA49rWxbWMUNyuNQQbcq8mTGsFkSqZk41zg/a6fQznWkY173
ZCbP3RtNka4ZSZwOXShEdropebnNfumD2HVortUgun4bdPpwW6/v1Cz0gfJsi5lc
1kMAPAKyEFiEFMAryQCdrDlDsBhMab143qLT8jVfovthwLORVRSDsf2VCR6LMVa2
GjtUFuGR/VpIYxTGMtbU420SO5+NA+ZVWTXWiPnImQfnzwRfYMVZyDQ0U9osmC5e
vY2MfoRIWV26NhL7RirSeUCgz9Q9LZvmzQ+Y2f6tHgW6BFBk2YcoIA8VgdxT3+tY
/RoOv2D5uZWM+c6L9JcESftLNQufZhWIwC8kzVJTwbefBuU/+s1QdUvSHgla+76k
nQ5ncZvp8cZVkt5j8pT1CawmK2vFAwaAEcB/nO2UfHKT4VoYNakiQ0cUp8ZPDkd7
Px5FocHM5IYeHTsi+YuFvX0iS14IsneV/CDjnrfmGeRwyFez/cGg1pN0oOYSSlkc
ZweOgztHxW+VKh7PhTBoLoRh/1E0rF19oc51sXh7RwB39hUZMNYpfjyz9g1XejcZ
mjJUD33vk+LAAwm71OImcqsBbmfjZdZkVIIH288DkZFNlgTB5jDLrXRlGgJvPNUi
NuG5zAbtMoXHnzaMKRVxkGFFNcQ7EuC9fKG5OEIai+3T+2VG0jbAnIdDsjLLqcPN
j1dMVmhd/7gMjCutYR8+QRE+85YYsXIKPzwIWC9fai1otCUiq81xT/LCY5dx90Q1
BYf2n+tTL56DoPN7hEF3RdAE8FrosoZVz/dn7go3/g4jkKspbIQjAJ6iQhsOx+eJ
yGYgVd2pvRSV5/84TRMJuU1msT/PvjIIxINq3vDAsIFIvIkiw6k/j39fAo/22C0S
CLQlKx7h7f9fFu/owsvBtkiUrO9exfCtmhSuN3W+jB2uoIP/phstdbGagxX98L6T
lPbmUBFt4BC00yEip1kaRl9NX3xtNJ/i8hvnZuoSEcnnjnljlbo+5m0xJRV3F1L0
2Qn3yb/Ur70YWVXwlKSTOn3ZGAOlyhDUYFPUZwIAXK+ALhBrl6WjjeuIxkGY9oPx
5WHHde+dctIJZorDIeOtRQ38z2dSDKwEUberF+UWJ+9R6s9AvrpP03+7NY8fIrWu
CyMcP+FxgJgpLBZDFAtEYkF3ZbWXplY75uYnkESWwiqPxOZY2cQ2yJA6RHenZISZ
aJmDTzWVzLUaJ9NGlqkKUavCYP/aRuWnsteygLqwvVZJxOQwphbXEiNvNwgMHtDw
yX4TAi/iL7J719F11IvKx0oDvJfGHbarBVntISc7vWDWQy1gm3KDwuc1vbWvc2iw
6VOty+EaCr99sRIZ92MtU/gyGtH3wwi1lDjthyAwThtBD+hggpywNPLnRsd4CUYI
FT52s7e48gR3JDhsKxoDpTCcAIvBj57PtevktZr1q5F9VV/ocyZDNelk44EnnfAJ
HelA2dck2AH7QF0pvSKfypkfoiZ2cL5u/qH2WMun12piCzJ3UTZIYVPFxOzQKWj4
5reglYue28A+Ux3Yl74zGeNaQwFjfnndq6QcPfAkFr2bj0yqspEXs+S+z7dHScm3
qoCevhpn2bVBgsIP7bREX2iCkoB+UTwLCm+HxfegTrcOcW+pH8noCvYA0VDkCIvI
qnKcR1jM5HxZkYFjuzpuxTYVip2kv3T+YHy/AiAksXiFlbzgzzZ/fNK93sC3Hs8s
grI+jHlvUbH5J91YeAx9fMQFFGe50020+Q4F68jRoQftDTEzJ9sbeOACRP9xmKAl
lcEr0jWCfkrNSAXYI8fs+2DyFXK6y6312vOrygyc+XOD3dqf/YGltl9aN1CrsdPf
X6gRnQ8my5XiZWQkqgMM3jbMihg0C2CMy9h7pM/r1DHCnTOeX5cGaZYHlAByhxnz
BCs2+HSYnpxxTK+z0licuOaYmrp1yX7paGP5VICaUU+TSvPPzD+9Fdy6Z8IEMvf/
ZN+bmWPrttecWbft/rr6rOykfkN+vBT94kqPhmPRwbvmrI/1CPpKP4266udycMOO
SXnfe4dL1P9ObxGcwLl/yZpL5OPMpuC+GxjCynWTD2qGcuDoJbub+vHDfk95/B3b
KgqV8uaoqK3SEkwZdtZuZrGBwr5KTWi5k6DeSSUtb8w9xfNmfssZ0MHMrrESnCOe
zRLySHQGypkh10xHWsG6MUa0nHBqCQ4/2KOsUQN2x58DNdUROxyKAf6wGWIhLHj7
Wu4b1XeKjUjmHpiaTY07/3FUPLKzT/gf/wIC+7lm9o5AyBD0m7lzDCdQv88zTz1k
xtv4+pJ8RbXdmbKZW04uu845vLB4gbgJduOYGF5z9081sQ06uJ++0aPoEFZl3Qtz
Ycr7neNbxJNENfRqwATE7ypPd4ACnBAnFL5Wq4QVAbJlw8Z/3uy/o4VQflP7D6eV
zOTUyqQ4wwX767GTyxGBBME88l2CISlJepZIi2Q/pmRArwRWVsyigIIKMl867tRD
iLFb9CJgWtr6xdxNwVOrBdDV5+PxyYBmd3JEF3zbbGW6EMKvSkr5y7QUnxF6UWrI
0mS1c3Btpn4Xbole6XCLPQ==
`pragma protect end_protected
