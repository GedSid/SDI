// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:35 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UDGdanVmE1zCl3rihgL9e7B629Espc+xtbtucuFJnBEM3eMh/WLiLi+zhMicTsuC
df7kfedHrFt+FQJSfl8j5szOiMNTQqjYm9g313Oe+0Y0ijNiosKhe2T0rKNZX4zv
z99S55Fd7vmphwHQTFdm852+hPEEyRUY2gq4t7iWlOM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18384)
1pagGJicQqs2GfMk+YHPrbTUYUcYf8+UrNPM9zgenVexeTu2Dke0MjHcEejRPMK0
5/2FvotskQhk38x0xSPhBBNOyUMvizx5WwoaQeDP2s8s73R9zeMQWrI+Ja4HOXuO
aBeWNzNzD/wY6lgFeaLdoXMlntkFDHbKrDX78SwHFoEYcXB8ZqL9ntu2wva9gp0P
S+GElo1km3Vo0a/a1rKdC3Q8B/wcuctkA0p4P/fI3Kh3/RXIApvfZ7L/5Mni2ogh
P8zzEbwJMSCPc3sDcEUE0ZrLSHSm23fx71a/0W0z2MxgbO9gayfdWzSXxXco7D20
xG9F7WMcagkevof6yRvRWU1NLAXvAcAnOVYPrFM6UQTsc+vuyrQA8IR8CzPN8KZ1
GFouG5CD2QhmO8Ldj9GZV4FDOOZxXZ/T+y4ZKP7XZRutlG58BklRMpMLmKijGqdc
JXEXxaNKIqkkb7ekXQ4RHPqs6WCj3B9uZQ0coSQBwkB4KjWtSW2Sgova22mLlhBk
duL/Shh0M6vTY4g4y7/UpVJUn+dVIcZuVLnvLI2QFWI9pHUQObBJp9jTFiv81kBB
23tumxFqv0JbZwLZz3XSBfpHkoejIbhxGlXV7ROe7b7PFSluCYAB5pghWq3vwNH8
HdkQEpAYffcE7Sy4cnSUeZWzLn6urbGPYRa/tUgzTcHOV82WZXUdD9hLdKc/grsK
5/QjCbqDiG91ExuMvMwXnIlBtsdCadCYA4Hm/6/t9E7hf7ETiYIbj2tCyQM5itsG
toUNH8mB1XurAdGjY5LZYFHcT0XXGzfCBGvLIA1Vyg7TScE/LnO+fYgz/p1pZsVc
/Sazh8I70IkTy7a15Nd9Sb45oQUkVRukE7IhFa50wbNjnXgTZqCzP4B2dB/Oucsp
9m6oQHbbqNx8TolJ2A/FuRkd2qztuHAAbr9w5SlRavnZR7v/jbPQfGFINoo4bQb9
Hlq0le6DwiDbze+U6x1r8Pl+6+IFVuZ1AJ+295yY7+RkJ9nWR++3Oo8tl6e0sWKW
/TG3ZcnbAhucYH0PNqhS5KQI/tluzhDM5DxegPmFjzEYCjLgpLz5ATrlzk1pqqGo
HsHlFXif0iNRIlPVw006PKMjZMj1OZhdyaMJ000cMcxK/dwTco088pXYioRVEjk4
jAoqhXPOY/7jdCT2xU5AqSQ27eeYzRhq66v1pHkTG9KU+zNRUcbHEhT1OBsmGHXz
lzwFXE1nVBLHl9e091hzCSTpmfvyuOs7rs0PGcSdichUgUhMg3dPGw5gTjktnPvW
UHL3VZSvB0GvofnxoocckxA42zHegcriqzndariPCl5wBKRk4Ct8dPjaL/gyhdxX
4ZLtTfwxOZ7hgimmhmvjyXekawDFMlmEPUIetwreMFEMAjMu0BExXWcWkuRX48L8
x75HTxo7YCf+gcA1g1lOmcE3Cg5w4DLA2kps4ID8OM0Y7KlNa/wuSsjj33z1zmKs
7uzy8Wc9Dv7Qzje7nPNrjHG09b0f4S+H+KY2afMjHuclqhmxnrSI1Vb7h02/Uq6q
skg+zip1lIsEW/utvDrQqCRPqLhpzZp1omHoPgaHMFCx79jmkjffxWUQVx+o23bi
4OYNEvwfxxTWM0XBuT3KQH0ZkaYszq6IbvIW0wweKia7MudhuDnwgxxHmg1TM5nE
Nj5/fPkJyZUj8bFm5uvHPhol4vIatTi7DCwIxcTmCk8rhuzQU6j+xcEhTpdHE/KH
VJcNsEzN1uzs5PWdFkxB739f3gDBSZGRkcBTJp//VnAV5U18eRg1UNFY2xggRWe3
vKlR/STmHuKX4pZMS9lBLtkUouvzvrduqquk75Ae3zQftBeLrtcQ+hmZkof5/HAQ
VbI/w69tgMpe2WE6UKFfR7cD7MwM2vYD/ZWrcx5z7WNoQ/v6EClVRb84UkXlYO7g
X0EBhk77jXb4W+0YJbj54owZYbACJndnMak9IgHLrzK46bzmYZfZIBDKK8tSYjBv
4dlbXQanpLNEDZS+Fcyx03gysv6I3DV5fRd/CynuO4IdpkgHM8a9zZVDRk+7w0Px
HtHXix1NY4aIMNZYGjd/ixkuomCx0bEgDcZAspR1GGsEN+unvoXaMnsONRjiZAgd
VXSODE4W2YiLFrntHF+IY9QmMnXk8UsvKuz7+9mFaINYfJoW9YAhzvaAXnmAv9Bl
rtfL/JSfOFMyPP9Mgkg6wA68dgmg/2v/aplyy7VZ2HCmb4kRGa72iUjvdqh9ssMB
Tqu2fuFe+3PuxxbScKSRSuF6kJRAJfx//FvMUC/9tHc5Ae0NJWWHYqSTGW8Wqcpl
0rzUIXikvhYFGKgKmsPrrUj7KGWFsAlZ62y7AbVlmdER1ll/RcyxszGwhoFjHBZr
eWEblfvC5wcZrbW+jaZqSo3vI6oiikBv7plzHATfGp3fz+y5Jc22UvvL37JFKJtz
vhW2CUdqWH7ICJSexUgBsOCfWvNKwBOYFnNgaXK1CwOM2Dw/9+ECFVERpP307yic
/gJwnQsnXZHWLl/dU3dfz9nNylYtAvCNB313WCODFPoOIq3SFwgbykvIL18ggO94
zbeFO/TJFNhzNW/IHpBU6Hss8hJrHTVdcxIiFt9UKdZW6Yze3iDcMDC2PHnelawv
XATtro5cepDoP/2HoIxziS6R6FHO4DDDzfLRWr+tiD+S3l+zHhce25NDjJZUnCU9
3LVYeVpAIp6RGt4cRnUfIuCkmm5CpFuRotN4cMWXXytI+7TUa8B1xiFQls46e79W
rYRaJRItGD0gm7oyF92LupXSI6i26riq7TN51gvkN3TMrOSNZZH1XMH7oQZGH1Ak
Xpe7srTz03syBcGK20dyeyvp9A74Ea/j/6/HThyY8fP0G60qLt5jB8dsVz/BlDVJ
sT4hz9wD8irh4KRuK52tzDv/fWlOcQu5HuzZ5scmML1Lgg1m8yQ8a5XmTAGru5l0
LmGzYwote7TFmyg0VBAKuN/mkJKdIjEm3LC1fthkknm+QmlZm2+RqvAMJLysS/sx
3ajqQKbrUC694bnG5uJKORjLZNl+AWSx36RBE7sEGDJPhgi1XTIuf8zFi0xaEc3P
SdGKVAJjYVgIk0P8aeGCKxrbehPdm3Iyz5y3qm1E1f+7a7slW5b1JTaVu8UNT/xP
qRkDFA18VQerUO45x96tnaS+OqyUppkr19JOp1s//y7A6Y6qbjF3onSaZbsBglwV
PeIkGZEo+lJn4X5882RrU0ff/SRdueHTSnjE0iCsQAD+EMbO/GwuQjazHdY6KVAT
Ivy7+uvD8hbWZcnkNNh8cVYWkuJNMtooOuBm1MHKP4rVIm5+9ZMg1Qv4ZwdYsRGw
0w99njIXv9IlwAcZnEkvtBRDYDSi2sVK5dho+DciNllrz2UjD5XN1Ju6rQEALDci
/vl0BMPlws15acmkydQdMuzewQptExbTjOM3dK15EgNSPRg/lQfXCu8DPCm0ZFLY
L3J4omZM8JYlT720ukQOgXyCjA01KWvucDN5S0iYoNvzsVgvlfyFv61S886J+/0x
nvZ4k8VWXIhcbtnnzSr+HDVLWGPp85d3KBgDaJm+L6jjF0LaBCPtqQtpdApFVQaV
ZZm8SHtPkmbeuFtNA+1CxEh5+IrxoWnoc7MxWCPt9DEBOTph99EfbpdxFd/9GqUO
JoeR8MHcu6e2VIJ36V8LhUXynscqxCN+2pUo5X4ngFFYbqM33DN/+G5AWwXRwgp4
3QS1e59jhayQryYm+N09VmBa+2hWZ5dbabx60S9FeVgRHHyWcW8FzZFvbsCegBd6
1qPi7Ch+WSGpoV1OWl2jIG7kfaSgJNv6vyjL2fMrEeC6+8DzyyRsyIyYQWSnoH9q
blaGY9gBmUo1zbKbQ8DtCL0hLgaWV4l+flnwGwSQ/ucSaZOT+KJOkurJnGlHEyJd
wBKAhzYz0jtG9ut3ypq3RjUmvdjtAEJ9DDZMAkidzsuNDhQP4lqHP0mDRlO7iWxg
0ffUQ8lQ2TOrn/nQ3fiQIBPCnieXWIhKAyo34mXZ6m7MzdlPk69dseyX3co3O1OP
sWQ5aOHS6TWVP+8LxYFhAjXh9kW98nNqvT2SldUko8su/PaEVyStQbWGihTpd16i
FtEhkGeD9ju7e+uNYjIMCJ81JBaIDF7LgxlMAwFm7mYjYq9O5BKjb+8g0R45LRry
cVWOGJ39S1IlsYj2VjjYuClryiOvAkNoOlhBXIcEbCWGDQmyV0UWXo6NBqPhMtDq
SFdPiw0PeLvfG2ZZBdwmDU9k0s3feuggzMWr+weT2pa65lM2s9JkIilUlLY/JeYb
ChnK5gcgeAxUgk9BuXxZkDvrXFnZHTXA8/sbDO6Gh2XocM6O3f9Yj2+Bdfd0zOEn
nGsQFOT8wYigv7pU/PJOy8eaSGpOq/gS29NzuBbQ4tNiBr7IXat9XsiAyWj7kKST
6wnHwZ1Q9VNBTqXz3jYqe9CC4d6kWFgGkpwmfM8NPEurfEH+Drx1CWJG6dhmdtK7
rrFpGgDIR5cuiy8CiaToAjkwPwTyAiHCigKiPJ9czj8OWRrxF0IdhZaKKefK3SNj
HHlL1fqwamMe18e5GyVbO44kufMa1FvXB+yBE4oUsqNKEd3/YDhwFLxKNMwRDvN/
tL8OP0hz2bvVlTTyWYYIsY/OCU0ZU0rJlfm6Q4oD+xiZOZaarATBD3+UxBFfJ5lJ
hIpbnwtVUz6hRfXV4pMLJeHYpwMrZv9XWxtcuSfJM/qwC6IaOeR8xcIPmrc4nEne
wAlf1gYNrUUpVmVrx43TnTSB/dCdQZR8mdGwLtP5NGb5HVjUJN3uoUN35pfiNGkT
W6cAOK6qQWceJK7ATchLKTlHvHkgJGR+kLZPSdi3OSvm556mRbdbhBC3HP4XTqTc
qzh726WMut0HnHhUrEna3Y+st9oGT9rvhVH2AOV32HR6R9km3UKN7httS7OsspGn
FcvKHkE/vb5iLP3rsrM9mKbeR0bIgiBr7stQoEhy2Qgr5cyjFn1FWj7rQVRE+JrO
Ffd0U3bPzJoidOi8UeUom6e8wW/YBx4ENe8lCMbo+RIt+lXELDA5hnskzPYhqiMz
sEOtZyl5+UB7fWAPEMLt/+0NZvO7627q6vTjQIWuTKrFAbZJa+dH+JqfRzPFA4uU
81mxFJPZLIYXZ2FGtaP3nz3uo4SQwyFIuVjCfX81uBl/M1G6/fE5mPH2blC6NlmT
YG+5NY2V3Y/A0Q92WDZARap7JGcLskA7SaohhWEftPg3/xSMGJBrSJmONYGvSeAm
dc/fWwBHaNfR6B3v8UAbZM/agOig6+qEFa8Y2m/8wU53oNBfiMdn6fyXEQ4cgOIF
WQEUw060Ne4Q2F/mHNgtVO8/NzBZfq5SXdwPdCd8/2w2JMsjrMaXT9PQyPquIxvJ
GvElxX+pXc0OZsnb9CScUNy5WfFsWEQzkZQvko3/AMxPEHnbgi80ic4e5xi3rVvO
NOSjbFirL2Zy/4IvCOnw+UajhA4QHEeNP//dFU/29lVgCmhJNbVD92dAseiLarx/
MxMq5DoESXRRKz9yea8KZnGy36QK4ZyfJsI7R5uihh5MZVGXpF39Xb2a+S6wPXQl
oV90VAHPjtyfGTXEtCZbiuWRtqz7PV8GjUn0Ut5E4JZJsyGB5qmzztYUwlqvOn9E
+rGsCbTSzK2Phd0i6E7PenuI5skJs+D2UI9gRiyeZ4SS3WkJ+8JAm+mumVtDB9dD
PIZYOBruVOdFnB4DfqkfCyFDOqXe7MBEwZvEOMiUNfpk7MtZ44Q4q9wiTM03sNdK
n+kN6O75YiC/oJC9D5W5HNms8bZsU9A4JobnXykqFtvjQBOokYznqHMVkqzXCqKH
Cy3X8K4NOu0p1tL0cu411pENDyYUJyPcX0OEdofp0MO0UECeboHPV0/vrLG6OWtP
kG5d4zQyxyJhNnZ4Vd9G0FQDaZ3wtTTQBQR9UykC3yOP8Z7fM+yMRnfS9ttwxpVJ
phvtYQZJE7KDmYpw97G/bQGuTKiOzF0PCBQA9pGA4bc2RwXNwWsthY/ff+7pIaaA
2P6psGd2hdEiACGwMmABXc9xhzdiKkU07Oj2QvN/Y/ka27/k8qS1dkMqOt1teQF7
cao42h08mWtqCI+v1yOZ6xKjCWvZYH26TqJZe3FwXGDp/OjYC7NEVcMNwdvwWs2L
mZQuKEzwnYeqPgVJTQ81lzbN+u7ijj5P4YsCurn+3Sw3BS003XJYsT1J0vkHlf7o
LupM3XFHbKFOjtI/ovaEjWMPY+Io6XiFs28G1rysT7s15/IZIFeK1d52lV8fl16T
zu/6+VJIwDaw5KGDfgQ1B/JYxIWU1wJkQBpMU99KLyfnO0c0hINkYan7N+IAYpiO
BBaivu8BsUP0mNdgQc58Q6gNzmYwDQMszjIpkh/gkuHQ+VwIYsJpTX4SCg6jWpGq
TtGJ0FNCn1F2X6X+qYbip0otenmHoKuhUCIxjebg5X8hH2vMNFNVHHcd7PH6qk9V
liO3AbrtBk13Syz2pWp5pyW7yt6nu/6DJSAwg8RrclLhqHH97jdx7OFM6PykBBs8
uUjo9bN/gdRAa8bz8ZYoPiMQyLep0v1TBQyVyq1yUPtkAhf3bfbWrNeu4vauhTYx
95LhTdiMzLq+kkAlamCKZvKWWG9TERGn7I+REfKrOrd95rUPNPW1F/6PyXOdPWYM
hoatYc5roddjJFXkgr1EFZdlS4tavZhQg6/vyZbpEvuHarcsATHjHHBG6F2q+ams
BN+JHGO5hVPfvuuZnfBLyemdctjZIRVmWVrEBp59vX0OwbwMDlTgY8crte4NFbmt
ZvPF6H6hipFfPxHKFU8w5gifoONaaqwxNp4mqU9s3rKmEPDzqVqUfIKurCIIVP4g
fZdJGEpJoBjzNtYc9oyrza6KDLnx0iKzQfz5jtMJ+1n57CS/bCwpptsOtej5LV8p
uv47kUz1EzLvd2Y2Nfm1sK1efw9DWouKOQI7JjS5e8XKVqrvTrIJ4L/2vPsLorPD
Gumju0K2SqFXZ63kAfqxBJZhc+HT+b0qIDCKHRuRwqKCR+IU4YpmGt+JH68eysic
17Q73GQegKFjzNtX6/bnPwMvKSNszq1c11b4DbR0BSVPugK84gRm/3KY2MSReNyC
TwyyoiQ4CEdnpmNhLITGdmpjCdm9oISXYooGlxhvb1gAtjRlMnHK4B+sdvFHaJoh
H11B2RcmdK7CEjk7IC7n+C+r7Ja2tAGJgq0cYrj73yWuvYgRpgxo4m1nDAAQCcm5
coBPpXeIKayWU+mp9xSlpaUIMI1mUjdQAV12xk7Y0pWgWZuYh2fIeJmdoa03Do5l
1wb3X1ePnbyDw6Nxe1aPv1DhwaYCC67tG8aqWaxyFh+aO5EzWuDOQgiDb/wE3IYA
WaBawaICn50JQxMy8jUqv+s8gOOmodQxwesgGrYCcSb509P0XXYqnwWiP3pVpb9B
t7Q/6IYeoRGev64Q4aQlcYjsZdoNTvF5ryGxIBL/6QnI4uFWuFsmKZ9Nq81Q98R8
KIOhFigEpN3OaDweA79kMAnkJjS5IcaroI0kknD3SNzVb/xs0NWTbf3t9wGCdfR1
IEgBdZsn6aQVrMDLRG50yAxewp77RlbIyuGNuTm+75leGc9ncZN8eAKomm0OnPiE
Jd6P1hv+njTA5ZS08gPdY+scpuCdE7an+4qMCWzqvxRKXuzv2yMTE2DB10wRN/nu
/oZ19IL6RZs89rljd1s+hFTS2/27n5+JIL1lTIeTqReBqidwmDtAK2OxEkfczrhM
7n5OFwwx4wSTN/jdwM8Ys6mgRWyCwOevXi/4vJ1/w5zk/N0Q9V68dzgyB9XaPR9b
UkTmw0cv9gFFYwS6FzECKIE5LodnFkf4h7Lv2XHXfD6EcgnwIfTp9Y188aosEM8b
Z6dp/HXfgyRLFzFiddb3KkpB2PMmPj5bo76raUWvb7wpED2AegPMOASbL1TStPhG
7Mstd0beuo+j7P9d1DCC6mZF/kYn2WHU0SRb5IUfg4JbTI9wRoFQUWejGseBF2Dx
WTIn0Og5aFYCEJei55Zsyl78H/cxXfOUgA96BXDfatrSq0dGzmR7zAMSiTNCZugZ
kpRvBDOjD/Kuh7IKiGKn/d5cExVe5i7ei6eciTu6woH5jkOEOAwFjEm0w8lHO4AN
gFCg+SyFcqc4+BCCMJOH2FonKL7cwXYFPyTt+EJf2eCIrsmvUHHSoZv7qs2VebVT
FhbIRDUhPZ8KE4AoKWatwgacyXGSXRO8KZjxB4+iqeqlU6x06HzBHb0SuwHk0C6/
yAtYwDsrD0RH7MGSfWoRuli0Ykbx8HhmXkQ/Tm784oVYM6sITdcliN+SNYaAY2aG
K/w9GMgeBIYp00/NiRME2lvOkFI79oDfvQfmMXOe+DgPArOZCEn3XsKCNnvA4efJ
MgbvC0yQaZCZGhOWlHWugaNRQsdOsssIMc4ih2F4vOsBad1okYuTNgGdNpvol9z+
g1hEsCNFukZ2VFSkWCGsr8k5EixHOex4tS4PI4Wtawkx+e1D3EmdJBGw2iSu+aE6
AMZNITSFkNcSRQOpfJUnv+XyWXaKLgUCEllenvbuQ+7qnvmxpORofmQTUG2MiDWv
arh2U7GX4ktDgzf2vsg4eAITRFF/+PBJHMXQMIs8fgLTLEIf3epwXdOX/gyF7Wt8
jJz1Ir7ldAE/fzdd8u7Lm4g/O5c9tophMtBgkeRpuH4Nd3E9cPbiEA6JY4fb0t0U
6+/4/BzcSA9gv4Ytpkv2oEfZnaGb9AaFFgDSmHg2pR/Mnvt1qKFDTRaZ08UKsWXP
fCqn9sFOJODDTT843dqeQkhAt2ggWM8qMJYTzelooroOjFH12xKgkvctDYagJb8I
IjFqV5dFT5OShZxHoithPC4gCc4XzKo2lc1euNJ7DsjMtKFmI+/cDv8mOMxptq7K
1pF40SUcSe8do9mxs7QA+vYYxmCjEpoeimBW65K8V5rFVi+NASqBTZF5TGNQfmju
t362Z1zQB7FuzR6hJgbaiNHTj0Xn+Y51yL8YfiI1rBL4OK6AT7UUca46QMTFVJa0
mYJz9numW12GU2mgLPv759NBjg1XXli+Zk7SFr//q8VWoyMm6qAgy7N+hoR+Dkge
UPPdEon8MacTA+SvTB7r9cjgDtBdUwFkwb6q862xOC0qTCZ9gWvHqWIhlgpGLd9k
j/anIaZUj9CeNe0RYk+zThnqarjLJMMT0sX4M0DLfjBrKP8Ur3gymppqwuv2pxlB
8cXkx41CnRvqXZP3177xfjvbshxUH+ZzRZyrZ3kKVePRNgGci7Qc1lqS2ygOCvl0
+HpV1hu/yxr4Gb7UrabmDpSoW93t0wQiEmiApN6u/++3PN/AjNtC6JIM+7kd1jpy
/M45ymv8W8k1WP2V8QLV+aieQwVfXcE4rKFOa8ntGavJJVdIfq8Afa0bK0oxh2UL
L9kOv7VN9ZIIQPV7XrMMpPqu83jiUP3kNHM/D5lgWD8XMn+quz4IO4Ul7D+HWTxP
UQ1dj+xJ51Fn/O+uWEtLJyE6cS6mY6qCmIkYauuLdR1y99/Gyd0pQEVByVGwc6B8
CcBCXOgK/A3yTAEUj2YRbRfl6D+biuUSkjoxFmyUEDKw9TD087Utq4tSgp2/CZRj
j8qP7ep4FOeIycqfxua30L+xBqQPmeWuaYLlUddi+bZRKyr3YL6v5+pnawxKZya2
vWe1/fB2m+FrZAQ0560hUR0IBIxs9nu8lfKGURIlA6wZp0qgaHRCAZlbjcz35Snb
eOV5lICYTCkRa3Vja/RL7udw/+x3QzFAqDpBmCcS8vgXtWdYpGMeojAHS7IFqiAe
J442QApGIccsaaHwSjoRMo+dTNjNyr2SaB5beAT6WDajnvFPLt/jI+SJxXJBHHLP
jhJLVf9j/1YOiyfoIu7J8KQXxMQ8+riUNbPdere9X6y0U2MISPy6nvycX3GqwuvY
ft2zjrgP2zrIbEIWTBP0DyRVVokpH0BqjRvgqJSUrEkWXw2Hs/jXhXYw+o8LiG1c
MKU9AFjb+UYECiKX3bKhKbBq3+oXeZy7ngYEi+SVcPjNuKsIoidMVBScOulcUdC4
8ZxdkEbrNTEt7rdbtSo9A8yNMDJmptQl88yu2a2lW/ws9H2y7hPCf9PM9pPHLiA4
w5Q/moiLyMDaRMwUyJybIPshnRz7prMQZyiaa7FrYB+PyS+nsnf2QAVyUzmymwpk
NmOC1FfWpyDsEfNG12EWAZgCSEhhlUYFTmzitRQ2FbjIPFgycWNsd/Wc1DVgQ+MD
R0qsWHLREkzM7nL5SY6cZX8G71NTHcGw8kGg0YXyNktXfXk1ioNeLKzh79FpgvCc
zUo9GYhVJ+C0gOIHsFsGxOrhw0IgsUM/kY1jYDasnIHJhGqWFQ6kMQvI0aZe2XQE
i3C/tTzw7hqg4mYhP5sAqB2q6zC0S/OE+7edRlT1n151j9yAYAhfRW439ZACtyeA
RSW84hZsYbXUDwGLqgH5IbEXCp+nQShMTJBaVavUl0K1OWqDT6GA6O3E6pi2nnpZ
KjuotXgDCT2PIpLZki6LkGmeYL02kxxAWthDJ+4e5iYbkTzd80FoGSivO+KM59Et
+YXKeulSOvUvhuQJBYhMaDx+X/rcugYTBAVS+6MhtSNx2dSgvw72+h8I4tJKv8++
KYQcpPNztM+B12zN31VyYdZ2jka1VjEGivBv7CQtqVcD9KnIfL7PYXwHK1/RS8wf
e18EF6TyQcJnhFXJVqsx1fDd2JMk+u1M8P78SCKH/c5pSqCi7aXdQHzQ+hKZLMpE
rgiVXw2gVLIlovQ+V+wjQTYlUonOesEiy3NO127VOVjmknYF9aJUPywSIR8hS6xo
Z/0uTtyTf4sQok7srv8LyqBGHBqFXdGYb18UuYmJ5Mm+A15Q0uAcrrCbfBepuQZo
/WrXMAXQEoE8lAq9jD3mBrDT3BENU6JsZPPYSBjlpb2FF8ICY4EAuItoloX5sExV
vLWIoSjZkg1k5zxfw5SpR1WY6ZrzRzEA6ijzd2+2bngD/hJwGfUvtAGmrPBvE13j
tfd8yQZHJfre/RxlGAFvIsFTjinKZmllIxXzg64UKkNA0LoEx0FKHqD96StDUq37
Mdo/oZYCxAmFk8Npp2784l430ex2Ch6nSd/uFV1rKTWSZ3EfSx7HT4lfIyoaEreS
A1cdabzsM1xXeUbRWmbmQ7EHzgTFKasX8cPZt/c2tYHEHe2kpgXcI55VeI6J/386
EK/HVOzHBSsokBxzQIlVsSXhzcdiLw1so0YymXzVRTVa25jR6aGQe1og0Oj+Ym+J
Vljg2EJcwvGYXJme9HEhnNWcagQnkVfCZo42TG1C2jnxwFY9acoPLGqr9aYatgSI
xUAkE1YdG44B6fu7fjWJE2d7KUlSkP0hBNCjckcQuRJgfs8U/0A42IpNC2WtJXqN
fHFkkeBiIPnTTk6eUg5wlB1Acz47lDhr5E7Ro7VMrJGoqxL5Dy6dypj1xTmuXxjc
A0OZJBPxi/Bs7mmsg0zhZE2S5zp5Q4awBJM9VMywb/DCHbu0o8rjurlOJPfKl3mB
bdlTVunOrIu6QQ9y1nLYCPj3CHZO/TaUVOPcN/RqouGjLjxvIZrFTy/LFqb3wKOK
i9TPkIVwk6y5k/jAWk94mZm03aP9snLUh6MjEZrRZNdSTMYlphazoZpvnloT1Nju
LO2UenlXunmTsAhvXld5KvUaYi21dO1zfSwM/M8+Vs5/nZFe3F6bWwjMaSXctFEX
efi8bsKaUVKs1pZhGL7n42OSXN/t4l5tqQNxl0VXYvcIfP1K5mGr1BUA+0P5TJXd
7aNskZaPcpEW8zrcBl7TMmMHOq8fDzJlCrJaNUSE8f4mfIK5svqMa64lIhemSTsM
bzKuT3Y3SBCRyOiBTI/aBXEYltUSYeCrK2RAYU4GNBqUDHfXcN2MBHUGU74gk7yy
proCmmXb7UJc6KssmIMylUf6uLTf0K67rNpu/Ss9ewSrJgDVOHtDTYkLwYPjgiDp
uZ4vAcB5/9Dr8kngUKD2VW8HZQx3aHqTn61XuLToO/2ON500tSak0JYQ5w7WqbJi
6neQnvbNRTcQ2QzWWWt8ByKXDsgBE1ur9hfTZUNBTDbMpV344qt4mrq0amIEo5HT
SBDUZc5dthyIDUEHm7kp53x9p7Kx9tKz1jBWUyYc0zSUVs7RHKUQ5bP4GvhxNL2Y
C95VmloZF72/uA2NERSAA5bkxHJ70V6lDCJE+iTucRxsb8Csw4IQWhoPhw9woqQ+
ZFuBzEiUx8/KLyJWRG5nfOrYFN36pbGeGP+vDHZkvpyN6wuhx6lBpK7n1ndnogXH
CgMYnIhjehmwxvnOnSOdFMwAMNcv0rmBMK3fghGUSfwHaJ7WMP0+SlB1/0h0xkNc
lgy6cnplD0/RglsVwaq+cPAL45QCLaXS1izLiG7vGAZIJtJrcpjW6wcZjxd8xGto
c8R0TXT5md3byLC1y2GcctjyABjW5acG4DC8nBFkThVp5iuz4yAFiEgpkeSCxnpk
N7+7jP3j8c6V6kdFf2646+kObfPnhdAMJ/BsdkXLjScG30ZHXxRDcI3q1S1P49gn
Uv56vzBXIeaC5K3ILcoHvPHCQsLqzxdYZDwx9uuphxyhAeJkwJhbQaVnNjEql9Zh
NQTnFdZF7dnluFz8w/54Q5R0JrN18i0UBLpAxh0Par4gW0AlVxPgpNn67bNAHziA
mZmgsbd2qzfY/29Q3t0HRM/c1rC8R092H+95HBlDNkL3br6ji7XCuVckV8cIyOOe
gCdKgmfdyIlc1NhDdo7a8ucQspZ3hbNXKY+NtJ7G3j8EXjSxC5Mu1WPopxqkRb1N
J+tSv4EGnc8fnh05q//o7T90dsWTYH6wniOVjGfpmOo0gdBJBNSjHK+V27bs84Dn
wdMJFdnnU99VoboSlvsru1MNFiS59kQgHlYStts+DHr1KI3ZH+aqG/Lwx6/+N4sO
SLK2V4isJWPqGvdSiAEJRuYVZAnMPaYR97dCP7h4XZO4mu3sG2jj6zo1enDgl8ZC
NGAC3tCXWXdurma/SPBkz+N4+YTU0BDnIkbv3FARzpInUDyEJ1yLzSsONNPP940l
vfIsUHsc57Ww5R1F10zoeWpwdu39+25P+0T5JA8kmS61xm9Ve/Ongew0sQi1CStq
Q9YNfdy7O+Kdb96imeZ2JiieMIl0k+OBdbiJqI41eTKjGAm+tSJddh8k0J88KgTr
35mqi53rSObfZd9OxV1EaufY83+wwHs0KBglHzLa9bFi3lvMbyGLg0L/04083Ccl
zsLXVzNdYkFcgrexgl8eSFHaVR+SXm/S7LL0rJV/f8sZ+8NUR9Fo5Bk73Tj1ov2/
H1Fv8Gli4RZ+JsZ4KRUm2WDqQS/yWGFB7qgH0VF+t3lNoZ2im3itB0pwRH69ha9U
EswGftsfsf5q6KaVo3xUCqbiAmodZnmbk0ztX+3uibEylyIhnfhhGiEb928XvHfQ
pamBdr9VXeUhjvxaa6teiNM4clViw2cjNN4lMmkqdmKRKFsNRWzsSVTtgatFTIoR
lzgKgNJjptGMGe49B9HtFiP1ur75EC5pBHxasJvc9bqBYZUgUVCUBbqtZYbFLrMb
/KjUCUip2dtkXVQ9QZdqcBCI0r4NKRzEsK3L8V7rSiLt0BwCaRcFifBKyiDesdDW
u52wl0oOT1mjaILdsmjftcX22cyI4YO9rXY1f23ku/aTQ2auRaFKXVNQMO0rZHO1
VCEb3InBk3KnxDv95BCIfEC4dTZhU+0afBF1uyhnv2z+jW5K44dDtTCBHPUiyLyv
beoBexpAm6DfJeUvl9DIjRQ2VPZNpxWv+vw/4efvz7/03KZ/mmoLr3KCE4GgUcJZ
fbqLm/6d4kujyPsc5/6WV2x6YF3TU4TdT8DWfWNcRYryr34nb79y7nfaVqGB4xNf
p7ZUcFKgAJ0dmrhIlx6/AqkEBdujvWWtISUmFo7GDf/27NCsJZHFjsipO+369wkM
0Lw8LnQb6uRrmlkt/QDvm4rWb9MBvKqJ+QThHBFIS7C47B6110Qx62JOYZVifjht
q443tSqerkJ0u7skRptSQWGfemLB70vxKOjfISZuN9Xwh5sXjGhxCx0HXx4MmlJG
YCfnaf34gVoIAG9N/zYxOJwo4j+HUCUhGhL36hysNhIvXsMewNbBXd2PL5eo186R
eQ7u5goOEssDSC8k2NEpXS/Jw7Zn43/CYL82mnO+ALNZlMEV8sE5kP+ZkfsBsEZP
q3ISdudCWOgZWY2lsYFj7hXlPM9I3fDYX3tJBRAVVJA5KTmCHqJsLNtnqMx8+0IZ
Z6KDwG26Z++2fyVq7qOml2c0IAVuu6Apvpky0rWsLVRe8vRRkzHqlps15Sz1w1SA
ja423HhW15y25eSZTDt/EgiobBDLiToszCirFFpTUIId3FCXInBneVlqEIX/Ga0m
okuoEwWFiX6qOfZk5Y8H7GkvlYxz9ornh1zsazor4AF1u11hMsBasF9vPnSRavyt
0E5rVHjxDOwE3hTze64Zg6qQRfNT3+8TT6PUx/rH/+pj6sbqnj5gFKA+2l9JIM2x
TQ6oTwJsQEBVKQ/MoWfCGnqG0Di3eB0jgRoDaSwNFlA9sibyjHovBAGCwH13Ohy3
Q4542zqPTbhueMYH3KaIHXMlx5xFVaw9PUIsuRTlsiu0iScvhtI5A+ICPfUhCnwd
eyUQ3WQX58h5POG8dSav2G7WITK02fYf5sMZOQGkxlaKSdtkMOxtWwKz+4hsoB/K
j7AVllHPB/79ZKlLuSMNCU1JXO6THivuyZidjX6qJlTpkeruBg05AHV75kBIyuGv
P2+3acZvfEP6nWtEFHX2FZ5m6O9TzB1Zm4ojnM/+/G0xOZbVrFVrGUDVRbazqirt
z988iDkGppHgnYLWREr31L6RnOY6HHmqTR3sK7xRCEOLDoNOwDLe4QKxZq8hibid
IkcWbAr7eYdw4vz/twnYoiL231rx+iyVBSjdTkn8oq6eQ7sdOhCTLjaKKhIDHoGi
F1KBXMVGmMz/3iig3E9wV1RyLxaE8yNGJ1n+0/c07iAtfGsCG4D9j0ccL3B26LsN
XYFplAqVRVXolgLa3pgSQhjOjxor/4lwxnLbv7ICwdV63FB9jNDn85/mmyULpJt7
v+gXAhMYPaWozJ3JYJgFJEbTU3+M/gvPZZsPxNRu51oD4rgRW27IU5AgEsheHhri
b0p1rwVUt4OV6Bro3vT0wuPT3h3xy3NYCIWS1VNyDLY+cQOBESJonHMt1B9ub2VW
fag+HQx653/fVDko+5ssyOn5pM+8XkIA+5GDa71jriWBW+XPchAqTg91xW5oW614
g+i1Y2Qru8QhJ8UDrEtUUVQiXF+4kMb1aAFRPuaOc+Wq9SUVxnT4kuI3kZi/0uDv
68iTNzZMUhXVVxgZ8/hNEvkhKGScCE/IMXxyp6IgB+00iQg5HwR7qIOWyiSxlDFM
3p7AE5xnb5oBMEboxRNz8huF9nS7SawqzpDcRErDf/FYVPazjgryesymta9/I00o
SER2Hc87UNX/z0waO2wKyHIF4tHXdtBMlr24449DikX20lLhutc3CuysK3rh1Bcj
8BiWBJL9LHaGSd3aB2+9zgwXAQG/ZaQFb82Rgm+SGWfPG7087DI/s+QvtEiZ+RGX
l2wsdu6hH0hh2Nzg36QYicrT+zBly0Pp3aHJxU26zv0c6QFJZCnLUfW+waOmXtxM
K38oaW5IEKKCI6j2NLt1kNtWzq6Hq3xo2HXEqPPMjHsIUgnugeOmxD2M6hJhOXFA
aClgrPz1bzL2D6zf9YrMf2wczpUJD1V0sqPTuZ0Uu9NdLa53CT3IlH2vgWc5OPGs
xODTpvy2xt8xhHGGRn8KLv3XGYF0gIq5Yhk76TXb8DKM/IiGW1AwDPFIBtxONPs0
Rg8VbxgAF+lgzBmWplf+FoLzyEEM0GN1hLhozlZyGIrkjm1WaNVEhOm1jN9OOLzo
a0D/AMG+Hjk8YQLZ9qmqrflfwSIBBlSm/Et68jf3d105jtvq5xHXhe1SkYcwz25P
t1+mdxMRVRXHJ73ug6MDDIfnc7kQFHKqcwriqCbktLRjtduW8FuavleATj3wrfZ5
ZCOGLum4Pt0P2EODV4CFdjFmTCdgS7GBQs/7IMd1IWGFRkU4A72I+UgjCsd25Pof
NielrGI9T/LX2l3PlobL80vYsnYRq67egzi7uAPe6EA8gfsDwS3eWlAeKM6jwWQ0
f33gy9cnTUQQKGnGuzKd7sZWhcOvbiq0qFCoKmV/yxTqhZEFw1G+1ZXYX7Mun+hP
l/InhnAyektEFCTOGmOllEQumLrv1hBrgfDXGPhWhSnHIXHJ/XBczYhHH+aUThvZ
uQbXeVtY56gLiEheIM3uo0jcpu5pyUKdLLgycVSzvi603RysRLratTzVimdOCoVQ
HhfVZBhqBee7XZNgrW9lxkKmTRs1tBFCmVciGgvZdZmwoucfwQev5ByN8ML0rUMZ
lpUo6zgEr9c9RRNJGS2ZA9iI2JuliZIQOk743p93I6V9c3v7eZ9LJdN35cpXruj4
54F7s+ua2nEw7vu0xrTEC1gavSICHL0Vu7kCHKFjTeILs6ZQ5nMtNij7gJVX4qXk
1SmE0ItAHKqU5nTHM9k+8TDXTlQF0zXNFRqZ2QENRWNcKHX2OiIwDehqz+whIxx0
tx8oXO0wmbtKUVY+t9kn1HPfkChu6xGfZ46aF5/ftaQxNOMttFyLmDXmPGZDvIV4
pVx1/yquzFZj/CioPilyQBGWrFV1S+rbM/WW7rnArg9xJ9WXNCE/lgaYPrI0Efwm
ym/12yTj+2y2cCNWMv/m6t/4J2PWVT1H8EbOs033W9H/VCEBS1h4naCLtl5N69ta
i8IP40DCnQ8BR/pLxh+DyxMIqj6TEvBhRaI4KGBT3jmQz0rcsEXywAFGGuQ0vM27
nMP/5Or0DQ8LrEKIirmtjXAIUFUXb8252LIFUEOYoGrm/jTjKjR3t42sqK3DP57X
aCfBGkf1pCx+Zov3d2ISBQyUF9qCKwCp2mxe8gmdhW0TkIqf6phSrcC7dDCdUvd2
OaLGI2GTfqv6wMn+wem7xazeM4pr/RReN07qNk2zpqthMY7s4fEL7vWmZf+6NLgX
PFwurczuraSXLv101SOFzphjr9BFiHfzJ43Y+QmTe07alwU3OUtPtSGIKWLtmfqw
V+lFWilOKrCpFTl6+p5i2phk7Bw77w5iGOX5khI0qEBeFN67eskTmD6zC6ligLBA
inmJTLQy67sKWvQA/84eyYio1XV/yWXlEkdrEUtMJl9YNCShIOwJoOqbJ8HFdbcj
JOuyRfeGJU+6c6OHkIWuB8eRRMNBufAsleGHkmrPK9+I4qOAgXYM1Y8+EW/uYUrX
716dJR1LvU8Fx/iAmBxv2jgc0quCLxd6VV3jGujg53HmDv+vwg5Yo+mt8gzWzU/6
C8+9X4iGI3plzUc3YAQnwNKxh6LL9/rACVZLTu0HceN5ROxFrlFTrCazLm8D4Lb3
6bpoBdv3bMX80RQ1gma/HgbnqYmQ/BG0Lr3g8hGw1lJGwd1tY0wl6BwGl8WJ2VmW
364s4vehJav1WfTakboXxXj1INu+pwHv0JOGZRmWuIew0Ln5HcSqd5gNhdCQEhod
7TZHfXZLZgz1aBDySypNOa1qfJL/7cfNd1iC26dtERIjuEjDjWE1Y4VK86vHNBOS
NwmbLQxceMjNvc735SKw80dwrOntqa+2ReZh1tc2s0QQWSorIN60XPrlI66P2n9i
/ogxABBbE7EHD8Sd9ZMCUe1Gks/PJUb87TGj7EtdhdOffYPmrB/gPx0ou91Ep5WJ
/zURJpYqSEkA9JvbTdDO8Vf1RKirRxV1gaFfl1T+KCQScdbkEisDIuGx9VwmN5D+
e3/iFuQOfA40B4v9cm6dIXXYGCPXXMm0nzBjywUE1NYeT4TWDWzHCSVbIfEotMqu
ZadOK47p/W3+KZhgHXzLuXlL8/ESKd2L1bHvBw/juKnqT54ML7h8Vy3fwwq5ewwj
p2wauoYzOKaORIftZ5NojmNBSoLMU3aC6IZE0uqsHiLOiS+G2LCgzzo/M8TIkOcD
37iXZI1RgwxLFmt/LgH9/U7abYKUqLo+iocLoHpJ3JqGAfKUDpoyLpNbqbIDC4pj
sudalaqdEoBqIFFfMZSG9a65XkMIrOU30ri2UuTOlgVU+AOkmq+VXfXTKRmADdyi
t71Hh9VjqhpO69ddfmE0Pyb4dzih9q2bApIYVdj6kP3gep9kt44mYJfK+kCWtzts
XbKwYErBdw1EEl+akLwJ3GsBFtSWOY8QUbkfyhJSSPods7gGWvz02Sk800ViC4V8
Nmfd2W//Kz5S2iA9mvkddmBFHX4ofngohNJ54AOk91+D3Q2jjStVUwrqEjtlkde7
b1rNDORZQMS5SnwB5vqNHGtqGNdnJibMrKaTD5A6xCY1Z5qwIc+CUBnTaeGmgiyF
AG38nCapbdmcED3P5YQBikA8s1qkzRslTkFnd3wTkBhVcKb4rYaklv7/h7ONnRpg
9JvNv5gmX6pcaTQomO1zO3iU1NAvKCBGr5vNccW4mqwPKOByLe1oFX2xxlQGUNsk
7ItW+ifsPaoA/DSUcv6ZFHaoR/uLV/xJs8r8jojBFN8ijkVSg43WGfuc1BanaJi9
UaRueG2am4oyn/g83kWhlHH6y0l8aTNFVvIDSHo9XrDMmAUtVQJZVjR1A4xhj5R8
GqkBnH48mJZgn5gd+rpaeWANIsfV23AKrQ8dyybwRvTyJUZPadxGBnq3/aiqIXFD
qMgA6CynQJ6lfQjHl5P9tBMkPkQ3MwfbD6j7DP38U6kzkfnUBM+knXpBhCwUGLmo
g/6NS3vMUk2A5FcHL/dvh6P9WzspvCx7FNCMkIOe6WFYAlXdBrWbbr2mi0r9/Gnd
TgxpUZqIqfJZXT/55wxvXAThS9N/uCyndw+3jGc4E/sYNkut6Zg1FUex57UECNCp
Giv+lu2yvP7DuLinoheU74MeT0Gb4hSHDbdfMz9hilCiZisReETiokLeBD4vGEaU
o/MrQ/BIUi+ioc1+uusudts00aIU4T8UG0VC/4/njtmJua8uHBNIktc8bEIh7LEQ
g2+Z1kwlcWci8hmhJixJhqU9w42DMYERNOZn0iGV+OhW8+R5VPtgfJZt2l3XJcI0
PgHApKrmlAZXNBfxkJUolq0SKMP5YRnGqDYTfW/DqB0/9ru/Kspvjb0lsYPqvi7u
+P0RBGXSWB/WeWlPs383qONMvT9ymbmIW89+mvI5hbi/fIrh2gTr4xKd1M7+cQer
5RlIsIfSOo+d/Sy7/bs0c9MeM5OCD4ctI9LUve7wszZZKwk+3PgVBVeKnzr4313c
3WlZvq7QY9+VUpWdJEqhrjaXyI5IVgY5L4s4ZVMrSHZBqhnl66uXJDdal/HOaEtb
aXnU7B7LYlhXa90SFk0bXR2ZGS4X3xfk+1SCG9dl4FVk9fmBh32FWyk9qjgiefyU
K45lnSAk9tTJ0V4c2kQhEr6Pfmw2YYfZxVMJkvMXfqhcOdhj3KMBtdVXnCyOTeQ9
C0Qfs8F5VzbcgjdsOW7J6WXzqP3izEcVhDQSIra3wUaxnKMZCOUY8eOOzbaXdqcC
xgOqUnMNRGwZmIYpAkr8W7Ilwd4nXNl5KJeDzjE1Fv7nw3sbBDhzmBrA9ZVLbymj
C+04R1Xllsf3H76GvFMTvyBNH/krsdmfLvYpyAm7QGSQg6iA/OrK5V7/Y2lkCEcy
A8dUB/UmoL25Cl3bV/aT+prOWesrlOmlNI7qI6lWtY+CG+YpXWlvYTKt4nv52EHJ
1ZAuiCzdUskIV7Eq9+icQGr1GToFcet0QzuDelqRP5/vZuRU3nemEPG0fqzbBUOl
LuCQEzYShV5pkyQeXg6K5TwI0qVCHi3h2vUFxwP8wXvNKwuSSRbdLc1zonqEy8+h
VjlFix+vwGfWXYD5zLdU8e4ZwvDR0B/+BAst6iyfRCLypOb26eHka6+1oBja0D+W
oUhmokhaUyVFjIS8NyHzp6n6rMiF852p/D/Oa2Hc2p5/6STdVIjyWCkjY7RmoddC
sAbzY29jxG7ucs/PH1pJEJwNImwlrDNtUePxz4Abp8xOZ3fJbvCJocFlcjngnaxz
ZPl5+fQHDJgkAQOnejk2du8choC8q0GhvqZhZ7SJ4PscxI8JfeRUequE60ESj0jU
hyO+358BfOOZCRVR7Y1b6Jxk8fpfj8dknYN/ToQXVRDyRDx6HQ7mJD/FlAc98Zr5
wxt0v5CADr9bv4o7NAH2u0fOhz8Irs5eCRewWkGx1fMg1GKSZAoJMCudJwvCLVCs
i+vhnWsUgcEy7lhFe0Zwb69QrMUNaqIB0Or/YgbEh200bK6lPWLkbSt52mKiUv9G
wLKM3+4t9IBU7CBG5b4ROGm0HepbYg2PeKC8wMgmi7E19lQwGjOJcKasLq9fRRcT
aRa31kpdHygi6FwGsQ/Abf0ERdVRGbNVJRC/NSEwwscow+5yqsR4CDc5mUpihaHY
HYP5ynxb60pZEVZn4tMJriBw6XuOdUofJ7IYNrVx5LPwsblt3yChK7Hq9LUCGK74
OCOTTNJF5gU6+UjFERyaTMqzfoHYG/Gh5qaaYPnDCenUJXqU+3KwnkgvNzaFc8N0
4zGtTtY5aPCsUBnRh/btbXssO22UFEXPnyWEIMjQETL3t9/OoB1cfe28gBC2Q+Zw
ymO/1mNMUshJpuWa9SyWsT688UJ9UJWjMEHEUnqc3XV4SXsihHkWPK+LVW620Cfs
NVjH7B/J7BvppbXU12N6psoq3B5V7tlLGC2lcpcFdaTdVZ/6XqyTpTuEzIVIWE6Y
LEefDspUXhHZl+QKgQ/odYZU9yq4v9ljnE5TKQExbSWB3/VIIjZWZPpYBNNHClB3
2l/QcUsCACthWR8BUwZRqx6MKcEUYLPJxjO11V60KVZkZ5pGW7AimbxLU6L4G66n
rhoe8kgaVUn7Wd5S21dDGciQGipT77G86GF1LqRci4/mC74aTNQ/RnWsrDwBDH2s
ZFtPwzJKaznyUxDpebQk0VWseGNa4r20chXtod83rmlq6CJ2EDRJ23OQ2S20uIrS
t740hEogxndKI4zZI5qW6j23PZ9qOGgG52KcK0LXXJjxKrZojO4cXo8cXWDJ/5Mh
mHJHsteI/zlnBJyw8cwcty50dop3d+Dhc7JwpOHzWDJIuAsiw1ThLA7d8G53OvKp
JE8Nu7AxfhKa1c+UwzShaqH4PIKTILUVpJAS4D9vbuv5buKgO8pVIoayYt/V/qQ5
Z97qedgM5dJZk9+7U8VQXxtPYLHcBUEQZWGSLwLf+yqodyP4rBB4s4bsTq0CC/SH
a/i/acjeYFdOtyuIn1luIzfuAC7PrXawWS2N9WbTVw9MBDt+Hi7vSlocFR4EgbHo
1X9Z/qOzzyY+u3EzIrpQg3pEPSOGe4KFdCOWOnI/fM9vHbhoPZchACzYretTEgzz
UshA/Htp9gulglMU1hLG8EBfr10TRJT6vVMoCJfN7H36keb4Ixjju0y3gxp6tfUA
rwq1sF5XbUbaszglTb5gOpyX10Q2DuANcLGLn3jLjhg7z0ByIObptZRF5ltjcetg
/ApaL5dEygScv1EdGg79Oh85CZZR2FWy0nhzQcjcSbexOKdIzVCbbr62jvg4m33B
rGvUOTGSbygD6p/TolDzll5UE2OCAJjn6ptFFUjwQgIQvmEoqvbAPsUmk9hnE7my
j993hJd7XVGtGhS/pxFTaofRHUM1mYAMFgX2QUdh27jYtFHJczfHcz/eFZ5Wkxlu
b3GKdortdRcR7v8pyLF3KVvejcWGHeaaTMOM67vBXcJ/s4yP7onXPmrDOBHEJhSF
fQV1OyFXehTfehCzX7veXGquyybEFUdEwz2rm81VbslKk6+9JvQ6g9CnJSTWAMRG
VGrnVlqbR5BsjSw4NFynZ/XuQk+aUKXBF6jI5Swzq8dpnKkuIPUlLdlyl3yXZwUS
qTJS8/Pf0oWRsUvsBMjDoz5qDJmVhRr4B4OY0mUmZXt64b+VfYS+27oFkwqVTUrY
MCclNzJ6iAL/UfwkB1RGI/KRHNzSy+WCj6950RHoGolgoImibsqZCtpQAYlIGvz2
8/yTJgqu1y4ft7ZW8ECs5InTGgFX5vSAw2x5KYW7ORZb4mha5ssbbG+Fs8SP2sOt
+iFv+oRMOXV66dD+hFSoL0lwNjp+mXV7Uqx6PXCDnXPh62s8amQ4C0N0GIyimZ7d
GVGIPwZbp+RxjJkXhXTqWE0mwXdT8eGX9N70DVCg036VNiJbZgKSIpgoUXge1GYn
khS186htcVKqBNVZroFrTWrPfLvYuiQp6ZUoTVH5YYUoHdgYuk7zoXc6J9wbn5zm
VJGJCHz4pPVwYbFis4UEjeL14CTYJ3l71SojIJ3V83xEPOn8AsZa4ThYR4uYwR+n
zeLZqDqPnSkFdOXCWbq3UauIGarCu0W+XUPf9B3UJ8dOGcNxVMH5MlxVmPlJ+r/X
vGbsVZaiWRh6XttBid7Sl1LOXiANS3EpElXa/y7umvxarnq1OKxkscexRYvkgVRD
8rnaOXBI+Nk00d6HF3auLnnQcx2dOBoNYafJzIu1E3ZiuZxD2rFF6JskcL1V3OTT
HfVF5ARQwSOp9w4DHoEHjtDFv84HdcK25j4ZofR6rYHddiY27xwCM40cGSnSyvpb
DR9DSu/Czx0aoek+ja1rq4C/Ojx7MpJbjg02MfNZ0fxAc7qLAc0XKQWa7Hg6GJJX
Gu9Ue68HyaoLUYzWhk3pMbLV/T3RKB0Nn3Z/n0u7CGtrd4MH1OoCtDFKg1ULLwxs
gcJli/HG8sXxFohLsL4XB4fXzPBxeraewz6AwsgfbRjCeZvLyYTT22rGPHtxaVJ4
8mHPq/GcO+Dpwdtxfd2H2sw+zAjwqX2chgjUvgtra3vFsTApNJq8dXTeKNwRY8ct
0hPguKY7PtKM4aYZarvaKi/+dyCN3H04/fEdEPUP/gHRo2pgT06R7NI4C/cVWmsX
9zygVUvEZb8Ah8iXkiF/hx9I56Q2ruUx6AlgxjLcQrb96l9XVtPd00mnr9vf5v0E
UDreDFLzE7bzk1xExVZejuigBlib+XQXEGedih6cd1IfwF5+/yO5RsWKIqDqVgsV
h4S+dj9mWAucMmvg47wnro7ch9DnWQViC5kGtkP0v3F1bEjXIMqc31+vAzMus6Bz
3bfWDdLytqn/IQA/lGLyuNMAtHRuUOVHT027MsSA90DCH5a3A90zOnPbsSRBGuyy
+ubSXk9A5Tuu03NMkE8efQ5GS6nFQ8ZClR41QSdY/lF339i8Icy/gXFrlrgMxQuH
RTR4wSZ9z3C9NcOImNSDCT5vIIa7W3Gq4vZA5ucCKy5/kkOH137b/DLHgiIvxjdr
FLMvAinF7Evi969w3R6p2cxoF07Otwr3xbjv+PbDI/qcoxd0jBjVDg4p8c6t71oG
xP4mcOc9oeUkXtly4W7lV3J9wmGX8TSZNmpkTDYAMPFZzEPgNVFkj+/zUeCnu4+m
AVubiWtq75/W3dWjIE23HuGZ0TX2KVxNqPT7A/EsMQLUGemqZHMjd2x1rjupUyCY
l8SA2sk7vvHaW15gy4zM5gkl+XSqqqO9m4trli3avRcloUP6bRuPpL6C+tkuZQJZ
bGKt3qA+dek9+p7gD+b2kBJVjsUcfS/Iafrh7BBEkEVVgedxq1t7OjbyJyA7Dz9W
jLihLM1bo/G9ndbWpWoRBL/ZesPx32+MG8ALOOmiH3v4eWOrrG5PAp2pb6YQl9O9
PkTkX+25X523s9QG9Zq9BeN/fPq0xoRb2M0aI4LAayjJ3yogOjGBjXGnj0rd/R91
i4hpFvVsGuxTT9tTe4QBb3XwPy/1Xzuf8KAeiiaav1ekQh3ofJwcO6KZ7Gyfen/B
enb5AU+0jyl1h/oI1LIHKz96WTz7cV1c3KPE9J4BzKqoUGAV1uhyW03en2cvOWWq
bo5TDFVG0oyqMYEOkvr8hKN+KziAXnHNt/qGN28RSVG2SFQjYZVJpdPlhSutPcbm
1AMkRRekMePTWPleG+58Cc4LSwcb/i0qv47hg6DiTwois4gI2TzTCdBeEsnUlDyQ
GWsJGcK2LfdCCIblYo5NP4mI0GuOXB0FJPXQQB8QINOx25N7iXFs7kg0EJZPUcEx
WO0kyqqmzRQ8SrJob2zA/WRiVRO3TLbLTumM7qAYbH2sG+eKoe3HajrRUsAghHMU
klToCKncWSicb31xgmwxuVrPsuphy3GMA0A7cfsIl6kw9jsxS4gbsMeeKcnRrR3N
zHrnINBKFQIbcCkk9U0PROZZh0D/47cWfRWDY7o2ibuxDeAG9XpB0D3J2c5Cs1Gi
HJpgRKhr0Xr208KnOfP1jFrD6fpaP4X3/VHh64apVl8g3AfuXQ6d11Cp3LOEM4Sy
orCMsQtjXCK6lpfxbmTve4GsUh2T+L7/wvKeREWRAnpN54ulyAQDR8olajYdzTdl
BAvxuq2J3T6KhDdu1VDNmA46bmrcddBP5If7f/CJNJNDAKTXNvse2SZ/8B5BK9Q/
`pragma protect end_protected
