// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:36 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VfJrCCPZVbnMgdK0RGGsbJAxKzc1cX8hpTtJIvGcKXx9rEXEw31CCWyKB5plvf0y
LIOurt+lyjSfI6iazu6b52o2qAfPYHCsbHzhsejJU3hYqArHlhlFQtT5yIk+COXM
IIuwx5DxcWnT04Xp6ZWRdsRb2ytM98NKedIdyUrRO9Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15696)
pjQ/OZMlmXPrjyJ03djow3dfJ18kFIzMK7DT8wyJSn2liEaMM3ztk+EYIit2nz0q
f3vjrMlyoqw4uI5XopLrji+4/Tr7jqmxKkonR6U1ERqQAJoXOtBdVwRJZXEJwbYN
Ew/nmQCwfUAbNw+iSUDzzAn9tgJRicLR8bGJ0cRcgxZPXD6MuqgGK0xjySZ8eX55
ALE9hfK8Qfdlo/DbVhVMM9+gud9OWZy1EMcUBwfEOBfoV+WUlBNYosoWuYAZjxCQ
KzEbJFnGGmP0Guc1mMsgYoPLUPvidxg0vMLbq2QwYJFURUsDWc6ZH8jAB6TiP5nT
s5B7TmVDBwMLyhSVWaWVQX7rlXTcSidBxtSWOkl6R12UasmtSZiIagCC8ZO6VBgN
SsilRI1haewzdN6SprSB1I8Zjkd5+1Z05s09iawA39b2lOAorMEAOmcjF6YGU1Ti
Q3f5Zo9E7deU20N/TVacPS/NHVV09VJu7BTIiJH7Yr8QVgkKnXQpm1tHJz+WeuYk
dLPrtIY9LOazKVwk/kRbDeP7PYjHqX0R/K0i6JRn/p1aLbJfpucMDpSCyaAHAXLj
WvIf7KzCPpA/vdr1NIvrsPp1w58yVHZjHs5Djuihkpa00cWPyxVYFYnpWAYR3PQR
mZG5veU10f+J71TJceAPmL3BjoKYkUapKT+8iQGeMiArjA/ZHSUJ5rpNnQGG8Crv
AiYj644NTmBj33hlsC4TcwmN1C/S2ntRlLVJbymdsQ1Bm3OZzXD+JudIACWoV4DV
Le7XDrydIDXG6Hb93APqwIux60oMNtKdZZkwLNpn3nPOsdT5PlnWxt3DlMJ8W9ID
wiIjRVJV28iKkasVSFXdGqukUDsphUMpIarpizfflO8HkkqDxUkvLS3TRet20qwk
yThIc7INNPG4cd986nYBudejMfUBnZRjbOGEFrr3bJoOWjcxWtD6ZXfpfyX76iCG
qrzPIsb5u0msgvb9ZMZpBdXkrpFidjWk3DBKNQ6yDeLA3llCVJSA5pqCgX9sc8v5
nXuuKGSZ+VMf4uR9mQWuBmESsdx8IpptUr245sSWGQcJHJ1C/+jgnqD0p9y9QvDF
GAvlvf6w/amMYc/+gKu5ZNvurU2dgym0CdVg3uKXhwlXr23N6wSWQAp9LSjTUElQ
xuurLmqo+ZTIEpeouogl1E0uMDkQjmqpxrp0n7ImjGVwF/dY1c7VgOTuqdyqc2Ty
FYc2u/0VOiRXP8d8q7zg+i9Erf7EBtsqpQ92Sv6fb2YrSJXc5xIL8E7+hV8xgt5Z
d4ag472BSCju2BJtnvvO6/fNKv7i78V5qkCxmV+8I6xOsUMXYMNeXWz2LgULIn0B
loEK5vBu4N9B7i1yobhoGGC8TjrXRJGEt7ZB8Wzfb5mcaKBcfClWb/ATSvChlKoo
TU/bAAXHLoVwApe4Z4OOQ7YiV4EySEEKjF2FkZMF7sLmD+nOpRK+PPrQr2IdayQ1
V9GFQAa/RoPxNtP2ZjEms41HkHetJGWrtf3IPodx9Dt08oDS7F10pP55rXwfTAHT
zMCUTejj7XPiPLAbSblyu/xsEMzf3sfkbUUyMsOz9Z+Wt2VRElYeTMWAR86bhjph
H9bxo/5zxqtF2tzRTMJezS7U9NfoLg7SIfa5Ih0cXJKzgWZnPs6iCIkMRay5RdVf
UhAfOP7i/Z0cK7+MS+ZCpevO5/ZIhG/Gt6cJnj5AXPCHC3p1rGl2yjCbNApdORxs
cKKkREt2pHKSXtNMzPTQyOnk4PwyPEw62L8uTMWslROdfBszSrMztT9Hnu74Gyru
hcbKAm4gLgdChP3Ar1VhRqsnf+p3g0WkuA9ZE0VRn1T6j1+Td8B813PTeFWJAR8K
p+9AVYQi6sSNZ5me9t/9TsmZdGWt7naDzq/4EDDBgX6RASlKlzZgoMqw3HAL52M2
+zovNCDsd8o55FY+mJatGumK+yy+SsaRSCetwnHdod1qLTJEB/UpWdTPCYV5zflz
88ACRMyvwD97LAr0SEFEQVQnRE1eDHqVxl3+iiLeK3ly4iqhQqOA7uTvZbM2T/5B
lnS28Wy4nltkFcHCSILyVipBZ1PXN2ah13VTgYXXF2WkirfL902UJ+APlTuXoYwO
e6V/ktx23QHQK9YbKjqspRWwwtuBHdG0TQj9Oo5wfGZSISyPJQSgN05b30R8nZjP
mQ643kbm9dkQNBPVM28DMuvVLnEQvP/J2HYWjb89ke5EZv2aydUWBqfhXQVMswQ+
yuRTBIzdvu8IS/p2UcsZiJXcAxRHKenXJk8iUjhyhnqqp/Dnd5jxdc+De01y6Fzw
t0xQe8E/SX6+rtAUb3iFX2WrB99YuqfIDkZLBAYfT13sddDlf8lWSfwMpRi28eYO
9G8ukRh4hmzAa6Hkyusymyt0BQT4eXau0WPPJXgkXIBwxP3IbxlOn+9c7z1csvCD
yIwfISVv1X2uamZEwUTugr0jI0ImLtEH+saaBuCtRXLcrNrFQfouem97cmwvZPe8
OA7DlsBuLEInIM7fI6FW5DuS11VRPnD8w0Suum50BMshnozxJN6VUGxcBI/hZeYr
Mnrg9JYVoToUoXvLeIiz3y1u6GMarJlJrzRiMgsQ0ZI+JTqObR+KhGnabcZACHRa
fKH+oQ0YmlfdSUFViSIpIaXkT410qxfSRU3F9C9cDlqaPrAifmBz9DQiaAa9xSD6
o4g+vjH8mlHo83YFP0hWpz11pqv1TQuMO9xDmuhHiHNkr4ATnzfVqbU2ULEegBmT
cFOktayuvS7A+VWaO0eESJU0f5efosLfRlUbmqK1oWlk+0nS6BZhpp3sCt4GWTYL
ks1sGy7CqOJBzZfUoA8iWy7Lh4S7ILYL1iSJs2MXDN/Rwks/SPwFUY5Z55rw/DP0
opXVFodR+CYWw0BeDRlkLBlRyYPeFsimfwYuI8E9ZXGuXDLRyOI3FEkKMoqvm7so
vbLY81lfaTno261hocQhIOugM7W1vXkSJaNbFWXeQ++KS6+X/HQGaveiuw7FEcIp
Il3jwkll5hR8nYUDEGk31etMhOTWfeN8YYP+YWYlXKToZinuLz95gLsvuRspBfmT
7H0eMNO2C0/MjPW7k7hnjTMCYFvmb2L/5cpDJ1oYo78eDf+aEzCqqOfcHThiI7b5
H1F/I+qvAZNjjA65gZgMv0zwitoT6/JYJ2S6lBTm6iyB82j6DYReP1JHO9IwcmeC
0ktqTffdUyJosAK42J/AvH7oo9qVOLH9GV/jBKSXWTmqy9gHoTSu7RjkJyAF5zx6
E3aB+J1LeqJzsV8HXHgrzTHVkwakTBkD7VGRLohPrfaNvaNtX6Xg5Qq0qmRBU9AM
s4BwkGEI8OPm4lxFefhXS/TSO5r3zy/FMWF2+jsmDL1Y4r4yWEzxPRNUMX17ned5
BfzngfQkiyy+zz+pgR9MFKhwhjxZtYNFtSMWICNjTSUIC8AXw0f3Pphp8ZQ3Evhg
alMVNyDlZ8xuac3KK+f84Lc0eruSm1nweEigBQvfNZVZGBgcdtupgqDJbG0WEqht
PmTfjCX5FzQ/8gD9rjcD3gen8sZMV1zQwjSBufWifz3UDzOJR3/dzz4BtAqwR1c7
15SUUNSFScRRbNFRs05Rtx8AAlOtpW5HTHM0umdsvm4UHDj+vYgSgUnNCF89BegL
n4moYcyjynnZH7YNDgWpiYrpkS6IghVWrILvmmdmCY3YAM3Pfb+eQkFQh4pl56tY
0SfIQiToy82S9LAeLIP8QBCfjRgHpP4KGVBJ6WuH1/Y+uWQS91utQx1n40hTrJB3
yvPqFf0CjTbNOKfcVTbWvXTOWgY0zPZv+BXxbreK6MsD26fLe4ffV/o3rIS8SVhG
qCa9ssg1XXgyulmGEDM51+lKa0l1RY3YIoH9odP47f1UVR7TUIAQzMMYaTvphTe3
WP/3/UOU3epLh+wswcKbIFCHQiT7HUietzIEj3SXKL4PhP5Qv0PkAKzCmYPQYRE3
wI3pPtLsdiMt+7GGEmz1CQHMDF5Lmqdnhh0WXw9hc0akFtDsZZxNXvH79fp4OCVJ
uxQRntuL5QPwckz8FpJxCVg8WFODMJa0cmfmnVtHpjtwBcFwYkB7J3dl8cts6WU0
XAuUrl3i3kRAedSoiw41fVG6+4gyhnpjmD/GVa4b9FpLcTWIinQFyttX1yBpjgXX
JotosoDrdTt/F/vb44arKacWo8zJzHrRpynBFRNDJI4DxGRyBDpGMFsN5qEscJ7j
GUIF5T0ZTWobOkG0vN7zMmya5p81QxoYUTzurNntWqcN2G+hmw+nwG4TgFy1p/kD
sSTKKxQKYS5M1etVjnvlwoBTlzKOy9X0dfP6htbc3yHtuiKZ/qT4D8OBxv+q6oyh
QCzBmjTbYCa/el3w4Mkh1pJadgyjWMKlZ/867O/HadxcW7qrpCcCXDDbUOy+m139
nSy4hgzhuXceBFwGrETmz08EAlEKIlbWTDtWFE9oMIuhLgipU4Q+qPspY1bCMTbu
Lt2Dl5afANWLb0A9wzIIZEePQ3KWwe9Ds33chUcaBhdO12kmgSZ/4Mu3e3QuCag9
/b13CyxZZy1DK35mQQoIqDZyPYmeE3rHM05nw/fr50UWr3JB6GbFutrqnVt4Vfrp
KmRJnPZfBjOFrvdhOK5aU6rIozb5nhJBW7xDOTYjD0XBjSw14SiQZAkgbwHDQsGY
MceXEIXCZnd3DGkcXzMXRRLVSAN40Vm9q03yNG4RoDbRBhk3E1zqKRMOlvsKyz6z
GGidOAUj3VSIU0ZcMzc9514MtL/jNAM/wnNo99u07M/HnM7wWhtMIWUt7rnjcq95
yaRc1TUvr6vqRh5C0/zpSdJP6dbaHP9dgMEe9MWM28TgP+FlN4ydvkE2HpO0GNbB
TuT6ZEtEWkgAQy9mTq5irgxHajBFsy0n6KiQuQEnEPVwqxyNBVY+mkjM1OkV43oO
5bF9xSp4Z5v1C0BiQXcIPnW9+faRZemQ4St22nVSNBF+C0CSUMmLm9zgGSSYsshb
kStrKR0dHutmXF3bNk8jd6mYIeLWkSgQgeaK9Fv9TPu+jPfLVBiIgrRUIKdege59
eCCPs4bcoLyBbDRZazrC8TZq16y03dNhfm34ywGvmzzHCCIBTjTRO7cVo9dB9IqB
8p0kxM5SRNiGLvoEA4/vUR7sdaZsYda/mx8vuBUsCsydHn176DoFtq3LnLKq4UqO
Nv2xCEdn5KXnkeLFu8sBIO3KQ32aI69iwTmytyUGf9vOOScpqnDuF6Bp0Q0Jgq0W
aaQiZ50115PxCBtRbdDv2Zpv7D73NoVgrfk68YOe84rHl4yKT17ir7VkF4iStR/v
BGZTDudY8Wxlzz/5WUgKMvgKHGSfEEBPCpFKLjab+xsv9av+0IOOmxiQ/YWbwfWG
Picgr2YGYpH09EE2QZEto98iVsLd5JfJka3ivNhw8jWSbdyWIJKAIk0Mb9o6p9KC
9x3zhNSg0o8mt9cdi0Tl6vBMHpdjKLzRlf2h/ZSNohxdEAWIVNw2Of/LiPo+kLgS
lYfN1i6cPC7JBgN0r5mPBHDMAdDMEQAc/1A0JRk23JAuwtHJ3aIna7VVVTJ3bToz
E3lJBp766z6AKGEVzl6aCTFBGes99kBQBr9uO4hVOayif1ihvj7F7Cx7J8kgCO3G
0CwBKlTIAOgUEC70uM/2Ms+dZ4HMW1xwdvR0mwRg7wnTPWXskeoYbOINUvaBMj/7
hI4WUvOOMnCzGC1big+q1+KgsnVItZeGaKS6ePGulyy9O62pnsUoDa6DXIzt7C96
44gvvYdOg3EfKQDRklg87HO0od1qu2xwoQPfoDS75OB20dc6eTDTca0P6luGeM76
uAGqZaL61auiDhoaNoCteMuRRORkRqNhWGcj72gziIpiZn6fzz/sfOtwvdJJA4OA
9OfcXCw2jPNx8UeXAJuD29oChohbE7PudO4cHAs2aHNn7UmAub/KYNWqyG8wDB+T
aynTmsZWTZCTHDYjYDJjQfEjuaqICHcv1sK02VJ6SUopUJ/L0pOmePnnYq9YoRIx
F05TxL9tQpMn54zaU41yy/m8aFmUQVGWX0LYIRlb6Vu/i7K9pUj69W81Z3G7a+ru
cR7+J5rV9FA4Xwd/xaH4B1G8uCE1lj0sP/Yy+FiXVQh7J6FkpoGQKiIQZj2z1AQV
KoBn7Dl6JmlEaOHO8ntmDzWGbmmvinqiinI2N4mhsMdmgNVr9KE3ySqE74u70vpQ
gXuphnRZvievRTQycIySfk2Vzr/M/5gIXPCYZPLr3Nt1kgX5D8axEYCJ4w6Niik7
9ifEt8HOGKjUhyAuTXWTidPool1DjIc1O228fdnDQvcA1CaJWzzsZ92NDzSOme/y
hEMj4LJycr/A4RzektnjmJ92FwiUQ6jtwooJsJkIJ0HRlXneCX8UaOO1gMWl5aHp
nxxox1YG/KGAvqcZ/bI791iyjIyg6a11V8CbbhOxWkzXUkDozM5cE0oSWvXtoB9W
T1PnJOPyae+tqDcbg90HVX2Q5xwU79zXVLRYsugm+Qk8/XYydUHQNiZpdBa0yIY/
311VLi5SoVVoaX1Y6Kd8kcsmvS+5ojURS7eJ/6f4vs7nFm9a98qABl89O4VyrNk9
aD2DeLDGl5Mk8MEeywW4GU/gZcL6E3O5mw0GksmUyQz2AdyMXXj6u9jgg8oR48E+
cuyhsCmEN4O04/DVJzyfFmIAS48zGm4gZQnuYyyf1FFo/NL6kAbX2U9G8zePXthE
npwNc9ujvD81CUBEcO/bUBWqQtz1QpXkL4M4Xt+pd4+cepjG8PmQRu1fXY8dbRvx
10cH4hnIkJx+HYwgYokjT2+SRVKFZXUZOtOCZeRXBONRz5gk5up6kWeyvy59Jl1v
rouDfW3bw9k4gHI3YT7vptO/1V+WnQrR+SWjQasz5zb0Gy9gB4MY0ptmIebMWdFh
f5tGkDKOg1RXRRbByuwZ8VypBFmuyg1yt4lpggLNnVDRWBZfIz1OmXFmCWYfGeFn
qViksO+OPHaEUh6Dmnp12tN63sviXRvLGMOGol+fkIz0iuLG8yfRy/o01mwC4wUF
yVniWjGQ+yaF8bFyI6/wU6xwhA4K/rXa4wRaOAg4YDSY6QY5pUCPhgUMWBfdTnEG
z5Ty7qNka9vM5efPkA/xlZU53L2dkmvCHP+SdHDcSNqCI1veLBYDexy5BVu5o++1
8Wem7b92N8Y629ExTZn0Lpf6uPf4ImkElfxiBpoKgw3ILTgahvedDkRC83c1L/QO
6TT8ujdVfz6eW/DaP6db3DaMThovrycsazahgoAOFcJG5Nzzsq4z1+uDsbkakwbL
ySX8tMVgJUe0q9xNwPv2DmUWpKEDJyCX7nZuB+Vw05xUoDEB5JzJpNhfxmwEgz3r
X5nXSjRt8bKoUgK04bU5zbBgFDBJwaK1nh2dYk8mGy48aufqOq3vuUSV9pgwd5z4
zBMzQ4eEOtiY9FxYLC68TZMz/vBXq951eP3cdT2F2zJkcBrGIN3sP5nV8xrUjxQF
tY7BgCbYx9nuz4C3+WqSl2FyAcoOhfDu3SZ4RiMLEB5HX6007vJ0wnIExoms8JXx
xw6vmjAUGN9cgRRjMe9ZuQE6zdz0F4QPCW4sKNuJNAbAbY2R6SyeIT4FjlCrIZkZ
xToEtvnG8hW8r+oFz81XJaEgCzmB0NrAopFyCzqWZXmxwU3CbdlOIAryalMgMR4s
hsUvlxBFdSKV7r8xlTstFOE/g92vUPTBEZ+8g2oWVQtHquh4w4NMrCkZ/rRAW/AL
58q1KDZmgXC1V5UfMZa1DaCiZFjj6d2sCA+5HPmNJOU7FL9lNlRh27vurOC+4D48
f6flBFbbKUTIiJbfFrv3kFvDoVifeZlZqx59BwD4AOWx0v+uj3E0xqvNsnI4GqCd
pGiglUQc9YXWXJ1qNA59tedzrfHsYaKEa6fe3a7mF0UwYtE5UGpnr8/qEvu9sG4A
HyOuP2j3wvBNuvs/LiiteH6kPoaM7sdz6CLQfcn5wqCpkAfMuDEOFoCsSRdYhrji
53V8jWQf/sVfBHIWqEnii63GiJApjcZP8dMNqmyLmlZ6zzOtG7alBeZivfXVtBy4
ULP3izIfgjttJeif1XDgvZXHeMc2vOc/opIxXUR8DaDuFvTGyg253N4bXbM6uVny
0Nmi62PuRUvrA2c3Eg3e9f0EylfED0xjjo1FNDQPD7HwNckhPRtnO4QOFsUCoTGq
1Xwcpv8tZR5Sg98WLLH9HQvyU0OfGN6vWbZjyM6S1LBau0unGE8vpXqS4BmTr/lC
Yjen6Kz7gMxpsQHyA+xZto+pmzFSdGAIdMn9AsOSW0l8/+U1I8b/zy4G0dBbwIvJ
dAcV2CWytc+XUHIGOrgA0BgpGyxwivLjYHy9NTLxpzoqYJjgDSAOhH0ID5X5qc85
5G0kuC7PULaW5t0jjmfSzZJeiOwX5W4NEgjQfd3K5b5UOUzCDMPcitjKasAyF4qN
YnxV7cQHi74vceX1k4arNvE6hl1+h1Q6LyDdudb1POODV/yy3u5YZ2vkYCrrbDo2
BSes8AI6YOVGNaSEclpiWPfCX26u3r2av1g3KuK79fK+AYAWRvRO9vO8o7+6ySXT
6JLwoOW2ygJGZOep6nzBiehDkQHpN1DwKZLeU7l4Ka6fHVkiN8ckFyLqw9AUgq7g
OdSP+gh1Wi8kc7wt2xnnAERHKAWmppOTPrgjnP0ABqY4KtUuD+V6uyFYN3dlL1vl
srhstPlUDiOeMZoQIRh8njzkUPqFJoUjtFV5z8tU5Wbgq/orBz53LwnWsxmSrIXH
ZWd8qAXaTvkmTp4qHcSKWAamK+1FWy+hYkLuGr3a3BXbhILADM7lXM4RSLDEFdIn
o3KkaEwY06XTwehnoolotsdfH2Ar8onn7h3mVQooeLuvFRig1N/ThurT+xKDB+BD
+nIWbDeXFDeAdfXal8d6xz7oJ/xZIYZDWwsvLjqFAODrKi/NamXE8h3kVPEh4rTY
ugphtTvxuulL1di1rY4MTQaTT0++Og/tjhtVjEahc8CvgxrmdXZ33tPu6QelnTR/
fD2xCXu2tojD8eUwEDTEcD6NZ6AXLRewxInn4wB5uMD8JFIkYz38WforGjbgJ8i+
mUd7Rz/4BTj+UWpyRKTmY3qa4DozqDqCoaZOFKqSkZllX0LQ5IbdbNouE3TsY/fv
+G5MRVnObhXbo5QZ2LGD/V5VHWfQhOjoy0e+7a7V1ZjePMWUQpIYZ1DSlDxto4wt
8rA4slCt9ac2GPgG9FuHFqhpPkKbS2BBkYymsqeWfBDVENZmTRB2NRoPV8KKZrgH
hePS5DwiMbkkI3Kqtdr7oaQWepibFiHkc2kELw8RHGqbPAWbK7JCuleuW2Vd1URl
ZYORie2niJKTwGP/+4YVN8Vuk/Ww20frRGoGlPlSZF4mVJfafKWu9IKnweh83E7e
u0D8yWPLM31CtPQHn1vjD9sVRExlOtiof+zwfANTGxED0uLihl7t3NlQkpqKteyu
lxdFhwwRjQzVCcQ7gE83ZWLXyp53aDqi4PHmk/DypYpfWZ+QezTsyKupBv8j/NfL
sv2DULQH8yEW6hIB7+NYRwzXdLTbLuliglAiFn7dauoo1bBmXIG6eWBfZiLA+Ij0
kSjCdtHLMrbgDBpXCXHjz4feJyqKpQuEaoVmjSKSyuaKJcqKXfa3L0bA+VUn/BP0
qbt63DaUjX/M8DQ4XbBIalG4FxTpIrltp2hSS8UnHefRE2+JnkhuAKYkd04RFZSv
xWeIpGutXoKoiQTkASN0eVpULXlalCphUEc9Pm2/gyQkdw+k/hIQl+09NHKlUV1W
wbdDUsdaggI98UoFT0QRktnRd4D7g94TfvbV6SPUIjrVztmR+Sv5R9pURW1N0Zhc
VZhE5H2f7Sme8mbWkXDdcGX20geTac6Fn38KpMnO9Sm+s7z3VmPjV5yJT+GFY2z8
h+4ODY5jjiHhoDCY7Mqbce9pJwBQ6aGsor8Jlcq+aI8DsoXJKmF0BxC+rMi5vcVT
MzZDPQZncaZJcZvj8JDYMGCmLQektnm6hdz7w9W3AmiOYTMtNB+L5xbJ8k7cRbz7
laIW/l3HEluW/u0h6ck02xhtH8Ymb1YwIlQ+G5QOkmBdVeVWi2Jm4V7yCYNmJmOE
8dd86CvGwFtCbmzJd+yPlAF0zjmTExGSsfPAnTom+BnY7K7tOQu0t+/Yj024OZ5S
cAlNYlzge1jETyVpFasVnY9o9xYR2WZ48bcye5vS89PZkfAddL7XjUvd7S94Docx
jUkiiUpnlDRLFSD/I3tvDuNdk8SF1RNWRpu3HMbGBFcbrbJ51aHM2RCEyWBQ1dsn
ym3c6qW1BSRcXho1i+6XUY7OSsw38TT0pZMAF/Gxnsz+e7NL1gIhbpTUtpxqO3iD
yPLVms3IpvaGUCNTHk2bxwRJ9+5PjqAGow8g/Kp0BLDin3L9fKSV9oKHKWX6qQkC
JXsCrOccQGNwJdpH9WWg2EDwC8SwSjZxQrN8nZZnTyk7PZKczKB/OglA9geUfqC+
oJOv1QYxYJ3txHUzHYkG3Xkd4s5B6L2J0ynNN6trNsLG/OuH1x9qjwoKSGqEqgXt
SEWcU3VPIGjUIi6QeQOqcJg9zUtNcOQ+8oNYxiPJnrSXZvzOq/bS3iSWE3Qqn8Xl
CQ6Ay/mBCTzeHWcwMVIZRUD+DTFGFtAvUbb60JqKwA4COZnEpIRbE2kzaqj7P7+S
P7LM8UDBNGfBZmdqwhg7Q4M3osoyPPU+duiO7w7JLnJXoeAMWktPbJfAY7YwRqaL
L+4sgB+tSAhhJ8umQpcKZ2TzyzmNiZd9dY5FxUEO+uLMsHxVKGUhtyDJIA9CLigY
pGyCYUCBHwQLNCVHNYp6+QX6KmOWsfJU0Mh62KkwUtPYDYDjDUG9WOTpuZTfsD6v
v/ed3PUm6TmmD8x/+7Svtirg73Tv4pUjXObslRswNV5fiMR2dgrEANeQWa3ti1av
JOLw5dRJm5XBHt6yo/DtbFs3tewUZ6h1D/XnQ+ZydAQWmKL5xjzaAWElDBJ2yAUx
xo/ctQDtmurHbo2Tjl200epLLJEWbw19y15fH6a2IcFTc8pnuZ2zAcy76x8rq7qU
a003v1c7ZH++snRxrG0Qh4y/CYYjTewCBHwL0lXMl9wXqBeP0oGK1zCyy60JqWl3
kwJqRXusagi+p9tSnljEdoc4xger/hjSLbHgqYlufx9PWyzDIMPPbZBye0whV5GB
SmFr6vFlO07y2klMe/vzo/MQoUuCmmZIRA3gvs/je+Lvwf51kwGRk7cXpXNotUW6
3kxmxq7JPTZJKh1I+wWi5p/oIDFTHr/wm+1mYpbI3hcoHTiwMb5X3g3tGdfqUqXm
eY9iaQhTS4gQaA+ZYFzPa/fprWCTLFkyFx0k07fFECjfDGBZZPf+o6qMXy2v6EGq
dn/zzLlDsB+AEogJqLxegTHmfmQbq96npzMGUMFaLLU5iHWrjs2ho8MRnQiA3kXA
/3+BMyQ8Ro9L1GDTnrOSHhzA9RnT1CoEHev2EakIrrURHi2E1gPfhHRcQH95BCK3
HEnPCF+XE0S/JjKg5kxK1DRHD+asGDsi47PDVY+yQPQHIpAGNOgBXfSDxrQwenPu
l5uOkhWltzdgoVuoTsuGyRVWgbMKIcPhfi3rft8DwapL6ncCiJPCP0Bk42e+iDiV
eQLmhTtHkC3q0aKN80tF6kOIwwOH8EQjiBgD+n4N1Zr4yUWREcqP7toL+OqUXM+A
NH1EWYsL+rzdFbtMEUSfJd9XBu89Amd5To4NHeEo3tvaFR6VY0e7e4caKXEuf4c7
d7gC7jW0ujAm+UcZTS+MNlVvmw8Fqu9LHaAkYyDQ/PMs1BKV3fuwZYwZlf8LPzjf
N+X42oIQkxCjhXqBNcOcdWxCuJrW9h7tKTyd34clC7mgRBW8qajhbqhLjviiB1Hl
FkujtjNXhJMqINzCv3AN4JjFAYYrAIRL7fQ56Cooa5tj2tcUFrJNdZv6ZgqMowny
VsoHPpL/kWZKlUlUCx9cJgK9OUZxLtbcDZRg2WjbTD3z2dOeJAZI6/PdsDRJmuyc
DsCpJpuX3S+o+HNMoC3lIdtvm7ltnRnuLhwp0vyJnTmiD8A1+EgsZlebB6/cY+2+
pZYgL56MM9/s5kGgPNrLMcAGWV+FD7npW/jQ6vyGy02JdNDtSfafwIocLBtwrKSn
4gso2VeMp1kC8YwjQ9sPi0v6POn6W2OI4uiu1F9PsggKLv3LNMFAEuUhFPpG5/lP
vhZx0+E2PKH4Xd7PED2QvFWodYpkk1jax1isv6u+ccN04cwfgFoevmQTyX8IYhch
6BhZQ0VHZ4WwCDHUV2KkHkW1IqWacCi+kNO4PH+v8dsrDEG8aadrPatndbq3Be3Q
JX7AhqOsz+Y8zadkBky6hh0Ay6ww2ICin3RfP4PKagUa1HmAl2mS5bMKA4kjHB4Q
kcPB3SQwDcUs+MkUsW0DoDgGMZ1orboR22Vqu69lozcUvaxialyK/jw9OOQ0XIFI
ExKC2uw4OqAp1ylkSLuXVx4SjzTvswBzp22khMqq+VwxMr5FoWgKAwqaE5QqQQKG
B9FHylnK6vl9Kn+Tu3CzG99dNu2XXp8huechj0b/KDMaWoK4Ljacf1ES0CmkMMrC
+o99sjHLGey/oGuVv1IV2CUCNY/QaZSlaMjuuTcqqPJMuqRLw8+W4FhlT1sF25HG
xBg7YKo6AEwQsH6xv2YgeY7Yx3R40fc+PBUzWaL+aDxvkJ6FpwdlSXpR36QqzK1N
Jm6sdQZdDtJIdmyeSi3ZaCd3m+kbJVufPcJCTVm4jTmhh2QGqOSFDDQnttefKoGM
SsDmWgZXQ4khOxqOEQWKLEJDYzWvOTdj7ozC7V8tvEJ4omLpyqHEua1POcMhvFdv
bOV8UenccP41DLfRNLdWIPhou6nHUjKuUjvTjgqL7c4wMSBYkcW7VgLXMuLn7kjM
rW0GWSuw7d8sEG4KzV+ckBxrHSddVQrTT0f0tQBeiplkUXOSx28HWCJEnhmCSxqp
rYqeBZTjnHPTRFdfoJeMwNfLFF0fflVx3l74PgxeNXSjBNb94nMm1k+E/hzl+FNE
1JAvbGQG6jtGhXN3I50VklqJpkp5omdXwH0uKB/nP5vI+5OtKmDNpwRJbsOtMbDw
BD3HiTc2ReQloGTa1taC7GPSkt8EU2Ltbif7bVJVDhc/GtAvM+KZI9foj1MYc6Z4
wQfZzwlJIL7r8/jghUnDFS0z/Fw7aAJSnq8JELqPjH+cLOMGglRZj8XXQdhPGuf6
hdqobmZNMfEmBrdMlTHsV4gwCxmrFa1sXUaae7gtMe0LF+qbe5badovGTYDA7iKd
z/XAIvCcqDPuoMs4Kt/TSi3vpFj0IoGxNJzo1wg8AO7MrnKrNvrqP/0QyHA0yxdZ
lOBoqCfLTy+hyZ1rVSydjQCk/Flug8Kmy4+/ItAW6NNGCoYj+ADAyBWscp86iQgf
3zC9fLUIrVtxusmsEqa9tta3zcca4mOoQH+y96xabJApiygEMnMkkIh8391M8TKb
OtmOfs+F7yExSMXle7xnE4NCgEsqrO1shcUJ1fcjSlWQhr4NT7j0P6ZP72x69ZiD
4tqS3VbvlHM0FXEH0J6eo4XxtUtIzAZBT9+JLYXdzRjtUeKusXDsnpYUasqZx8jz
OE9+yuDD04SXnfup2Ie35J0TqOZaSJ038BZaJ/8reDWTx9FxNKRH8UubrTsja8OE
K7Cb1jvkzRDRYQsE8O51+uX0AbFSlTYHm9NoJy9RJ8q6ZTgmkt4D+R3A2wdvpcFz
gPjPifBErDYbBnr3XrE1jokrGbbxx0AjZ0rcoOksAKi7cyiGfj+J/p6U8iab+GNq
W0RLFziFKS3L8OXMqKvbICXc0/JtKZwe9sIU3tiJZiCAePeW/gnZAiS9a4caCnIm
A3YyO47LaJUkbiJJnPlRbtzeXR7MITjpD5k+tISE/WAmuhkJ3FYIp+yKRZnuTY1g
dxJVxOM4D3i4HcbERNiE5kYQUsrulThLRv1vEpp8NV5LXwHDgoPlGJw3/xYJEUeA
ijvarGA3DqLk3i1vekE8VpSD+OUU1pzvmvUSMld6l55QJOo4RArA+I1V3Hwq5qED
YnvvjTOOgfWGK3+65YtmnU42/svdPV2yTD55JMhKcwiWU3Gu2aHaYovzgSgdo9Ra
3iYDNdHXH218MmXGPYTBqfLFKXyLe+5pMQkgYnINGChSOREzZrwXXgp8prvwsGam
QrpRWXUhD67PCbZ5afzfy3WKGievNEzQG1ihQ5gZOOjyRNlAmds3uW6tDZsDW+qw
bJPZ45TimQv1ym0ukxecZu3jKnv+cgNmWxm6rht+HzQJjZiJytz/s5bN387MfYcd
VaQyzSHhx32lfoqsGl73NJFud8eerGqsnqi18N9XHf5UvywzWmz4N717gyKzYa4S
cIaNDnyE8S8VGd2L4bEfvK0WuV3HHAAbI8Y+KZXNMviNrfNVvE/+5aXZMZsGSLT5
0pONYKo7kyeTXzggvO2k8FyUwvwDkppFm12T4f1agFwcetMbQqxkfgfco35/V+/8
8Bu1qSvFR5ohVHwiLh8VucR3H0XjegoHDmpsWgWa5arOAKkXDYz0pF0DJSewSB/t
krCZ9qxnwtLpPdipFwD6fNOpME6gKKQfxwM+/GSWhttLClej8ThF9lZt8axP6Vry
7LyLiVJAN7XL3kg4l0VPCF7cTPpvGB1kv4um/Y3joEiTRSfzsTE2y4FD6oQhmWgE
k5dX5WhYSEZXQtJ9VE7mQOVTrx7v7r+z9wO0CM5+zgcBUai2X1uPtHydZXTeNJC4
pVhWhex2ZEGAj1PVfuFBtEyPmu6qAmoaraH45QPr49q6/Wt8xp9ik1/RFJUb/0Eg
DUrtDP2vmtShyZ4lHc6ej/1FF2xj/yKaYHMeuSSwsxrBUcB9SDh8uv7AlR2ra7aM
6lUZIQeppI5ld7DXiBkPveR/NZ4nPeEDNvr3oI/M5Cz8JAiqtU6MHYo3JP3EEUS0
z9vlI6Pllx94Awxu266QWbRRzivH5biB1MilPJEEPSCYrnW8tXSdZnb8Kb+Zwd4U
LfDUl03xG5sl4Y0UhimOjVad9tjTAjhY3lZvtDpinSCejPouZxidV6Tfc1QPpxAC
2mQQlr7g+9WXsbCEvZg2tAAB+TTxTvGO9kJZgLsv3qGezixP04dWZ/s71vGBD7HG
cT4V1EnPyYQoQI15hYfIZdIdkPu/WesDvVGNK4iJLM41tfRoc3rcNQ/JS7s2z7WU
9fYuT6k7UeYo14PZvHoztv3c+8f5dlvG6eEQ4gw4UTQCIven5nkzDxPtDy0iTmkY
uL2spNG8IppCgeiq6O3ryZhuK2iI59uOFu4NM5pRghnrSx8VK/0bIxITs5Gcfura
C//qQ/vTmYz/5MhOrgvdbutV2fYTik6GScVsEEAOGPmHnAjLtld7BwnEKvEP9KlM
/MiujOhbm45QqmbBETlKdfUZKF9q1Bm8AtOfbEIbyZlH0wHibKpc3kqUjrOQWpKo
vNpQTUluOM923lDDIdHqWu2vGgmO5Lr/q0UTNm+fjdiMeBM7YgOXA8kEfFqd/x2s
nkL3e3IM7TqPSiLOsYb08lolQ2NuXmboqrKCIUw2MwkuMY/zj3KxmM/lT+hBjwwM
FeVAF1AyPM21TBobqmyq5AFbkFGAst7r74fYAQU8rOvLGg2egfaUwGYfu8q5ZQF+
QbbUrnW/79HP8yoSmdxEWVn+/uHWQGUewmg3Q/2nPbRKX4BjePlhmit2swQbOcqI
45eRMf928AfBmVbvulj3BZ9bT4uNF1yN8DmVpOLZpgdazRHZL3z/uPxDKBsEKfDA
BMJxyzw84ssOP9pqVHO3WTpftlHSgrPaZ+iWIZkW8xzNTjBPkSgFht7mgfo7Ij+J
wBttWRv3bNyHupgXvD/vvHEES1AGzaq4h/7uIawEt7Q0Hn4xdUyfecd9wuZ58Onk
AtDeLkdiBZ8+gn1g/YmkXmpHI7rDMo6EJAQq+TvzHwlKN8ZShp0jYtVICVjDOzum
oMnLDBimXzVaDPc7I/L2CVHkK0FVqeM60TbTTUm0KMVV8RjIVdc4QTdt/HQDyPW6
7Alge++xvCRmBUkYWrCIMPgg1y9w23awIzsR048vuEkST2oecDI5UaBKEosVZCO5
zfb9hTaIhrAPx9aXBLiBHqIFBGs83m7QpIbInMU7nL8l0aVbeMj94nYnwr2hTBlj
ieXdr34bjGll3oVZ+tCL5GN4K+QKp47tzYn1wDJIMtb9NGHvFJAzZNpW4vR+FOsv
fTQupx8Vo6VfqJ3WtGUqGtztFjc4qbGBm5HcLFVKv8GNCEe2PPvD8R8j2DLIAoRT
9tt9lyfxGFTkJZ2nZEUCjJnQO/coCSKgBvhXn3TorJdl4ZPMXQjMOwuqZoN69Qqz
z4O/wb+BYQ3oS9eMvEackL4bC6EqDzsTZ2uPYT+abqQ3bLMq8RZvYrxH/Mf60wuU
PWNpxOTKyhIcD6AXqTvoSyGesXuhrm0hOgkFNr25tSFg/dS+qHstuCPbMTdSOjSr
YFoCLkJhJFCjJPG5h0Jdl4slhvEJ/p6JmnBnBqo0WvBfZLiqR05o7j7FCvePzmeF
XuGkO5DD3qZbRvQKiELtQoY0Kx9rkzFjojfqnT/3kqFs+40jV4C4M4onakIbf21j
0Mskkp64BCmHRQexadhpCdGGknAr7KwabzYQFOFBBFn/HHAt5iqKF6Mzuj6u+rHR
cTXVJmgMInIIZ6yM7r2I2MOuXT4crjNeqnSA/o0pKwlSYsxKK/IyscHKilktzCIi
nYTjfsK7TacVnv5OKwHotKICbG9NU16J8/BQbUUaW/jdtyMAJg0igM7WecU8ut9t
ONWLAjWv0imehmupNYxb2u7k3YKa0u4VZU2WIPqXvUd0zTo5yCBa1UIwjUMbB8rm
ek95k0tvmJ/1xSY9p2SJWuZBZ+/+Dd0Dcw+FqeAQeB+Tkphkh8Yk09TelhKVciV+
1NcERjXvyf0zBoh+BFMXVz+h88x/ysxsPo/1sauTdHbrdmohSTQCG+TLgvNn+s1O
R097o9AuJA9b4eOUSGf1qO14nPzctZ5oqwwE9jiK9eCMVpn2PYFvaErgL1vSHSs0
PsiHYToIWvh7Y+mRPkdtu8xeB5yvUFmKGDkvqzxpK4OH/JY12k8wXPhI0FdzZUED
b94POovbBwucawRuYxX5LY2JryYdSf30yfI9Pmmhr1cYo3VYAx7vQa+CSkz0lA8C
YdMgOeqUIC0ntbxUnbkQcSEMasgPGczIAz4EX/q9s8+FDv8lgnJJr/FtsPxivJyc
z+4zYWCYM683tiManCONJ9WmYYOFGWPoijgoPoWmBEMNipnODiMY0rz4UrhA7D5v
NsKhecVvmM6C7gUv02Gc7o7vmINXmxrpooKjE2hVU8gwOw+Sx+xE4z2yF9vwEeDX
8WSb+kUlVvS1wMVEouho/9eJJNZsfRjH7rhXxQlQDIid0+G8b6mu1SvjToZEqMWC
O2wXQ8XFhJKCjZzwWUZ32wAX1iMAfTcp7YqHbAN5B7fbGL4RaI3xRKrsc8Ih8rUz
L2WC2rnmNO8T3iO2UWwzUTO3BZDhd6MUgyUxVJALkE1O+x1ErSQfrnfl8Gtu3Rsl
fmCD3GzuhqBBENNiHSruo8GFIJKvlPib82pKCUbPY7/vI0sd1lTIZKVL80dm2e5k
aIZpD67DgQkZCmAi5Wq3nb+zBBIi93UokXTXAStCH3vLuxudLD4V8+Oi/acoRTjH
roYmn/2wjgqgadlpBMsz8kt/S18XqHXpKkdKl7g/9ruX1Qq/fVicATHlUOTV5BIw
mxd65gq2tI5b/qbrwhxM29aU9j2+ZWzVu7/nTUVfFC42pmnlXaH/ZUFNLFnfneka
VqBkgk3wsVlhJzQFulSTXtTUyAYZGQRco7jE4xGD+lHU9Eixjl9QPW47tds5JhU2
pxB/rAx+4WX0cKqoBhRA9YCchaXYAOuXBKOtdhjqTUUX0M0ufZuPrh43gHaANTAV
JOy4cY4lxlwnvq64jb4gIQqe58RjoAY1293UbUt23Wmh/Zze5IGptN/L8geN9lCL
BcKJZ0kot4tpfTrHSq7UeddWd3QxMMFoTHNNGJVxl6Ggbttk/2Qz9QeS6BhqzIp9
eCL2LPy7VVPC8pv8h2142ZxWF7xrkDUg5BAqt0t4OiLOrGJtfwhLlMnnAWo5yaWN
bOBS31WuiKIF8IO6FbGQMRTdX/hAwpdalTfqqFbC2JMfLOWTAjqUu5dsN3gvTAxK
jfSECi7Oe/QeX9YW0V+HFJwhATymcvGBRsz7oGq68rzoEKwe55vAjY+IM2R/Zusv
EdzxPMa5QPV7iEnsV/Oj1QLeMu2bCpY5xTLvjY1malyCSJjVEgv8AOQm92u8hj1r
0snQUORmCwtFpZUEqqzmmWCx7H3V+/BUj3Q2iEXATXbPWvboSL9NFtro/lKy+ml+
MwFAZX/WdpCFU+qJ41cOUyOCDOmMwOsiwYh1iVQWW+g1FGFMJ4EzK1OqLwbrRAFd
8mssydCLnizN3zPH4C7OpvsgnvlXY9N1ObRPasbhdHprcJtVqQiPo4vMLyE+WKYd
YoFt6JGclV37lh0q246EuPWzSi5XLw2/i3/FfBkDzvUQW4qMXO5mFRj4N/+lw5oi
byRaIV+zqbV+ee5PJYvFYnlyVrF1uPvfsx1ZQx178KRdxZKnq/nEqLB4updQ7Qwz
sTAbMQMrHGeAtvB/sttrar9NfYya/IJweifvtfIDnqruZ95FN+EwYLVTZUsDFOPb
SQUFh3MqpW7E+G6sDizDyx3wEZFds8+4QiIjc4yv1ophyu2qSh4+QJlIYerWMXH9
XtT3+zW127/2Y8EZbgvF0pmScSbSRdBija5AZTQBG3iBgPflmlagWrQ7nTcmlMn+
1rhqgOABPl8TvMMBBmfnMbR2eojVn0/2EX1yMmdaPm7fACel+AhmnyD8U12W8cBH
BuJWp3wumvFxPMl0c2ETMjV5a2+q2DM70Bz75rNSxZ596w8+yi/ntOXQnRz80C0V
PW7ZoRpTJKy0LD1eV/glzBhWQL3nfBKEPcWu8Ydp2evzhaiR9CwB/WZU3kGCm27T
d8AxVl7Naz4L6C8M1wnT6z3RaGSNGn82LaazFseMrrK/m6eN6TE2Rceg6wbflC5q
uaJvruUMv8A1MaGdergKzRSi62bp6K3t4R5FjQJs64QAEBTiWm1epGCZVPTFsu/z
lfiyCUTbJCZSyp8VzmW9+saZocjmyTDWJXU0B4IIhvmH8MR+AL9zho3bLDEfRCy/
TPkQmgg+2Kq1dJFDcARlgEHyj3GOwZ5msOX1xYyCpy7vquSfvKMB6JvgO929JLDk
+IRS8Vf/ydNXLpeear+2U4uvflViNWE4TM4mVW5H06S3oAoCBViHP7cuUNZV9a6e
z2TFEEl90o61oDZkClk38vjwvYmY8ElgWz7YjAHJAeCXv//CydTDfoD9DFWgq6U5
hCqHXRBv1+/2DbqmIoR0Kr7ThGthUxa+inpNzwZwXd/XWUp+TX/s8fXp/sNtrT3p
9s2aZ1BMgkdc0os3cBqvLcskDcIDoo45Y2fgo+gL2f6c7kX7uMOVve7VEUo8Ts57
2mUF4YY+76rKpcPYjT2Dx0NS6RfFwbsi/cQhXDuyJSAHOdvBF6mfsdK60lerE3Kf
4IfMzcHmw4yHfcZSszq4MWyS1TErIjnCIRkxkTL0JGWdxVnlMVRJNv9NhE4fzKRd
53VgXjwY5Ubu49szR4XPctL6ZiWnBd7gE635dXGK0NBncJutSsCXJde1cDJBkziK
55eaRGTZ/bfH3Me6HuH+Rw84mYp0cSvlM8/o9pHPhl3j8Tp2uVHFKxcFlo3ihEwb
/4+ISIATiRNKo5MRQ1kevqELLduguZ6Ah1+OXDtODQCQjCKoOaXd35JHa62R3irT
ysEQDNOWd110+caBF0jsgGh7JtRSYqaoNZRMSYe/6Ts/uP/EF++Xip4Xe5ohGKNm
ogQR6kqV7K4mIVFgSB5GMcA80RIRNcEqXK32i1N2mLkrfPSIjl9xppW/4n1stRRW
Q2WoU1JNvJXEaIvLwJiT4CuYONouUYMk6KY8twPOuhJQANhQao9gZ2PHunzJVXUH
yobkeLW6SN8riClGte1r01ov/P3cJQQgrL0gEAkgWBuc6yd1wXqARZmXqTJ1NYXa
3k915NdbndFg79Qj2cJwadA6pBh1QrMA1C5xiPZUIVKm2fHK3FuGu4WwpU+8t0I3
W2FSCxXqqR20z+hnvIgw2C2gFi4J7BuKIVCuM8CUA3T+BPxCpXZmlZQSmDp62o2e
x5ObiK8NoQt7QvyfoIxSBDUnp6po3ikVPOPqIRDSND+LXG4FujzsKMp48qGRKUsk
QcuUf+Yu4gMlk+mAeQk7u7IxjTasS27Zl4seTGDgVBUSuIq6iAEWgBc+ocu3Ikc4
YIwQymlFHUp6fOJx2FBP8ZhVnrVu1nwYEWwckgBbGLVlY6JMOoKNw5ZoClyHkYAh
2seVH+k2URbFFDfaOxvm3V8LQjeVo7/X6qCfMP8i6J0gI19WkOJ4V7sPcwuWlYP9
KqS4cXeXe7nXQCZS81dKTV2RGFdxWoiU4WNGDljqRh8pGWRLNN4GxFm0Q5mC0A+u
5zS9qfgJoAqwx6EYW5vsohu3lT9Qsm7sGm4u0lfKrw9f5mtnPzrHw7rvp6d6CD9M
7W1za7LWG6A16jKvg68omVU3oogtYbT27nE8yVS5jjm2ww29VhSpKLLp6oWOdv1M
OMrdAUbiL2oB3aj6KtFRCukiVPxjJHd+sBBSlBJ3BBbvOjTqY9GWuSseDb8uM6It
UFzhBzDDfo319+hF2YmadJC3uM/2M1LsGBYAaa+XRjJZva+zPWo4tAJmLkqxYmcM
b5pH1l9Ht4G2imOF1a4Gjq6JgoVe4TA7BqfzdJy3+CPBLd1Wjhp9LvXKI12G8Hfq
`pragma protect end_protected
