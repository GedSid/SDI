// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:39 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FWO8NqUoixzPkxkTgr0KW1CNjsAgCuszFmgrjy6YTrYVjWL80gletQJv8i2Fz+8H
MvfC4O2+1eoapHK6lwBF4rwkUGUzjen3Cm5q3S+GVbQhSs+GxlXYA2IZJOXTfaqu
8wO+8DsusyQw209VLxPZac/uDYrnNIDvD6hlog3vMAE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13344)
IY4LvTrmqBwyrmTNUGHQrRuJWpzcoBZdeNsodGkDtbK9QS6ShyoRx0fxLTQr5vgR
OZ88f3mrAhYhSBcAOTBXrDtbBLjjXgt1tH8tla2zUMvujC8m+Ax+wzN5cQaKYKbq
rptvAAQeamEYDl9b61xzCEYZCpdr1c4Gf5+Rful0rjnzneTU+0AznTUw/QulYo2H
Oxfski+xtcmdAHY1clJ1VMziJQkyfhHDiS+6JltIePSdT7ebTQuFH/SSvT3XJb1s
4xuhV3S5MmVum8a24qzbNNOHzPckGLmFRSq5fXHHvmJcytXIVUKNY8Gk8xX0Twed
TI33YrcEM1bWRLOqFFyAlyi8kJYaoqPXNX3O/9Ezvz+TX6dLMge9nHRKM9Pwuzc7
xNDDLlZLoKfllkX3so5O6RXpHwuAUouXGhjKaZbnxY/wx9S7fTk28pgCGBrPw9fD
yNxUyTtLffBXscxpPFSNCaCQm5GW9SAtnVTcR+CJB9pxlzbYyfmJJ9m2daa6fRTh
AFL9Gv+2AnAtNFulIlvP91U4GyqmazcoT6Ja7RanLvqCDIBzuvWJYFKtTyOkQhXJ
wGPt+ZmzOOgOChKY1a6dPgExpYSFHlxPbtIA6G/HdlxkGYnI1MFhjUht0N7fE8Xt
LC0LWiMMvBl04YJx15izfdqc7w1ao9RkVHssxIM3V4fi+ZNQkrMvYiIIT+SRO/2P
0L7AKszAhl3Umg2ta6fWJJz4X2Ok7hSDTEiPIwMtP3z7jBMNtGJcZrFPeaZ7iLss
KdLRI9kFowJjJmEuAwb4vO5e3Xf2vBck0UWwz5ePo7w8AUfMHHKDjePZal5BH72s
N/rOzn0vZ9kG8aRSf83KqA8c5cMhT4Hnzya5koqsbGekOTjDCARFXdFtHcboIpti
nGnJONcOO8qkNCBIkvZP7YNt34ih6SSWItA8Ix4oN69f/60RWtHKNfnxygj0Ww0U
GrAZZEzh0llI0lwUopSH95i7zI5l5kCYalA0PU7vXPnP9iVaaZQyk6E0LiXwDVef
MAmQ9n3XKhCV8XpQ2wEL0+jJ4IuFVNksrRIc8uYGXZVOP7L9pfEdmYo+0HyTNkjV
juSCDMLWwcEaXamySeDZ9hgx0wIVf1TKAg1VDJb0HKgWgP8rUBQCX73sRKGF0DxR
g1NCm59armifXtwyMgoNzhHdFwebtao66Ep9QQo01KfMqF7GamjOwL80PaHlXthS
+HHUgbKBOdjxY59o3uzvWREYPxig4+twXh6pqMfW6sE05ZLYRCrlk7404T/TOkTr
noDaXryy0Lh2T3JvynRL8P1s8xLoHtSoHR2Fwv7dDGjDeM5R1+rZTX51z6TOfPXh
YyT6erGYm2ca3GifNoWYwbEUM2rEoRvEM5BLFifn8mqeCGgapQkDoIg/flXeoIaF
yIX17WrFBcJY3PfiL1tTgyZj8IJEVNEmLRKCFKu2oms2Og0WNpflOMy8IH3zcxBF
dkOZ5wgt37pvHxXJuP/ZIVsfMraKMnSxtK9ETHt8WBE6Ftj8kqcNF4Iht8s28YNi
ulZlI/xO+YAitXCNmvnb56H5JqhGTqlomIb31hEc13HHOF6E5OiKU03WBbTQh1lb
GqInxvUYHcDyZ4DC4bXHKLhpeHJmXXy5QHZWO8JxxS3ZMWJpnTY//XGqJ6WhPuva
lFhprwbcyGzee0mNOAWJBwBh9Ex4Qn8vzuGr3LapeQ+Y5JdZspMRBSXx+Vhwav6R
kpBGLXVVr4xfxzqHFhjcQYfT9cwcuvsy9WmnxrK+3aJNadV0SlQmqm5UiYZFtShq
zpunC5mSR17ZDbf1Ijs25Kt/B/pmwSxTvJ6jSUsOvT1YaAJ7d54GlWCh8iN2uzjV
go3jukect6dEir2bV4Wc+S10ErnFDZYsVWU8JuE1e86LU254REJ9pcYLi1z33wud
wvnhLa22nRLgIM2eR8QJvu2zT/R7DLnp/8P7asgU24AWofLXZZUEtK/E71DvQwWW
DxgxwRC79ezJJ2EWd9tHMzH2+voXIuewqSpIRIAvhjTkqhILP0s1pssL7hVC0DG5
Mz3+yHAulPDIVpcLW1YXZkNTC4QB5TFeb9KJxSZz0gEqgfXrysElDBBtxXafkDrZ
48gaEA8Q506XKiOMDQnF+yE9ixxgCxauSJ4JNAHGbFsvzQQB4PkFQufbCsSfJHY7
YkYSlYh26+flizGn1mnmHZUAYtDfSdNQh87t2e1rJAmgmIMA31ijmA3TkTpngOjt
SR69KeaC6lfVQ8DuLRPCsxOkdEnuZQHM1edke/zkGo6osTV07/OP/P7fSLa8tU9g
TH06EqeGmGC0ZUCSkyxDXHXVatgGlB6q8kfT1qWL7MVe8PaW9ECdr56M6ejv68RJ
YKSGSMykOq9vlRsdc26S3zUj7kBRGa6dUG0nVgy79lzcJUHI5lha+WjbhBm5J+3t
3TzglwlQkox9Fkx2Psk6AsOuaC6ThBSHgeJ3dzIFHxr/4sLb71+oYWqAv5tY1zmF
/Wu8IMslTMOvM8ddUMpaf0GylDIuhafMm3QKa9FVp61QnchHisgaozWoxgcxOreU
1bIxvOL+NvKPJMrbaVjhRAJ+1RdwZIwLt0sOM02XVekChbGPRglDCw1NvdAZMHp6
cJpk9/bUrCqBos8eDQXBagnHozmBcDz0NgJjucBi18nP3utckcTO0C4dALt5No0l
porKl2U4juTa6DFhOFlaxAQ20N7ttush2Toyg7Q/qMVkvnDmPJ2ncGJsitx7tzQs
Rur6d4vyQVoFNnRo4oloVyzW6R5cy48dgpRpCQr6vsoxuB7D3FFWSuz9DwMEwcyg
fwrvh3e/9D93gG8qcA74nFCllo9bkdDOudxjUax0xLuzkmbY205T4X1+HuySsOTv
P7iuzuLXtb42cqGvQjJwZSGJTB0x3Mh4sw2DOdfbOnK1g6clPjTqdRfDAYU2ZArx
nzbIQ9CeQK/jRD5ZOkamwk9zM0RWLt89WOlTkUvyIF2lcoQwaFZH92dmfSp6fsEW
xUP2uKji0OSr33xsEeOltrk3TgplmDaZC3pgznBAqRUFZIUygJEIab6biRi9g+oU
wdmA7NmKcwJGdlH26bv+PYZeM3ZU1wAw1kpFNB2HNb455hRKhEKVTOrJn57mdf7P
FdQ/UIs1lu8A+8Sm3ft8nMOuUhm5V50C77z+rgGixo2Z85rz1eZaEkaC2BiJKAzG
T0JxVvGNeQ/TJCcPsRPcwma8xvDNCu9TGvCOcpiWbDK8/3O31a/3a+Jp3FE7o4NE
xqagTdzSLecqun7Q9wczsBC8HeB3SkfqMoBtQnLa9LXV8Hcmw6lVbve9QFyEJAXH
1DfICPwcFfRthXL+lFED4DpRkhycsYKbfWrQFXpGEsTD70JZKbVSJZYQW7sJ7MCe
CZOxrpPCn88rR8bZSq6xjmJ7vuWbnG+6Y6I8qyUY5GgsSZErBSslINjdI/bzMDWG
X4KPO+6Tte9Oxgg7g5ZoSM8sP4QOQhJ9JVfHRRrEydUXKKWm8ZAD8b5Su6B3ZYr8
7CppxGLTb4bsmO6ydUDYCKbPyB39PAXNTYnENLAAWfN+Da0bVsf5E6Q6nmFllJZv
SEx6K6EswML3tErZph6Kcy35zJGpwxsO96w7TAaueRkVyrRxp51YTn9NPZ0l2S0a
+guRY5T7PS+36zD4UCWfcm2Y6ZMWgRKoeFRiWs2AO3xdHNRzSntEZcb1wc5cX8ux
7spxxmQhx0aR6XS3Qy2GaXnCKvhEzgFENnxn/cgNvolez5UjCC0KxC1louUtpHLF
+8+SAfmjItHfFm8YZsvKodNNz2qinVaO97xkX5yFRSR0zVzR86tc+r3/FLzAf/TJ
tPa5bqWGuKQA07A38HZHzgzdm3T1goUrdWmT6N4lFTWWeY1ZuthPu2VleBZpyiJ6
pV5vIjY0Eq1btOqVO/cQ1iItl2fAo/w7UNO45zF9EYf4Me2cJrbHXMWmbgS3vO3Z
PmoheE4wp2BlsrMcUVSRDyJz7xI7kynkEFiK3fNsSxmzcUY+AvikaBKrRlTXDbWa
P3URziLiZktCE7zj1kFJUsTYWk/wkNTGFsMMBgNDsAQclZPc7q033oQ0TpArWneY
2NhfMEBUH8NmBrkCP8q/b6/kJYV0LxYVggcY0t62g2LC14ZUYYnaUsV21/8xFFTn
eHAxkw8T2k6vq8TZpJojQ/FO1BCfJMr6kXmPevsrv2RO3toBFRJRI40tMt+Cr50h
at8qRI8Sval8FrLbkJd9QONutqgUjgiY55jMgLr9BRPzIOBwq9cv8EvhZ4z96RD9
/P6dm4uSWZPglR5OF2y4xv0DA0bLTIBDRz3w1zikXQO7snL65XbGDbyYW0MKnB0R
/XXBGNYI1l6+0Bt5on1jbiBT3FpxRqL1r1Gk8NvkLwzIcg75bP6SBGEO8f3d9C9Z
torvqlbzF0Tki0jpFwUAO+FrUvaNCORq07KOnv9Fv2xr5MDNT73WUmafxuHc48TM
ea65Of+bLxYO0NEZE2D7bNmhfbj2LyP1E44VWUdZ6Oj/8B1NSh6ak6kJTAqJaVhF
RJIJ0YrIzQ3nd+wEDtzfV51n9/gFWqia0VtHy0o85rpTk2ou0NBIotBoehligJbi
a3Nc8tXmYSgSNTUvKjvEtvMZJSvnYVhTKSs+op4CiIgvy+xiXdRWguljF1eztx01
/lSsyBdsz2UWVOwrQVI4JQC90mVsTMM7Kh8RnMOQ+fpeUp4c1iOwZjWM5wnJU8ru
vA2pt+uOb0XBNbG6vqP82v5Vwffqsq5DwsEaKzyh0mnpeeChDv1ElJNriuc2Fclt
ajtUCuT43XugiYlX6eAp150GLclDY9PCPEKIw72eMVTPJlwWAtiS8MdEUrCxIeb9
/GXYWihcBHNlI/Kwd+9+a5uTFqGJ5pgzQai0DTw8YupS0DvgmEfJl9NtEov16S53
voWPID0oleNLFgqRvaEbVG4NTPy+ohUFNVSZkUMLVJ0s3M1NVqQixbj2azfYLQt6
BHkf62wNEhmmRxWQ/CT9wAFrwFOa7Tk3hllsFTaXtfmsT/L4fwbHZ1lfWmKfBEEq
L5ZqLPGPgOQ21I/IS86y7ePMnLx/AT7QxMFXDgk853jR8XxbIlQkqCejFGDFgQ28
fvSpAx1ZwN7MfcxmYrWudZB4n1eGQmNvUyyfV3s2sBICHpgPNdrJQHQMtnAw5CZU
ZSF3/UinJrwutTVVnlc4hcqrNcB6hH+1bNPXsDzxCimCI6TnD3lGeevsbLeuQBLV
/vRPiVZJL+eO3GiTL0XAf9CmlxXv864krKmYtyvxCK/Nli4B8Fz4iVqxncYVrhHv
N+wd2YkIZ4VW37El1FUB6LQZpSph4qVo+tuA3/d157vELZRJUKJKVW41MgJPpdkU
jBiUE250xbbdHUZPVglaUUJAO2v/dlwQh5RKABnVO6HrQWCXtL124bf30F0eMwul
+dsUg9jSAYRMfSdAGhSBVAYDh+deW49L31XVUcYzGP7rwzuUWKo7LKgFAXLY+onL
GUOfXlfZ5oFw2AMuU4yWOzYwWU/6Wf0tqdZWueECUjE0dlKtEcDkS7VCa53miI+X
CQgW7B4WsIjVlgWiPxp3KpCpyN6FSouLGoozWdyErBCKzIrYKXBqgbqJIauJCB/S
xpA0a5Q0GysCvRxbBQ6jfdlTUMC8CI9HLEmLyqB9JORRgy1HStkohbOZdWFdToRk
qHTxvpDyP42nrbslpb7eoiu35PebWYauTJLKisulIyV+LM1qwzr1Aj/S3hUilgM+
3yGtvB7rTQ6nQCI6IeHjGBZ3TQZa/H+wBubFF46wYA+5xZo50VrJJg/WIGBIHpaJ
xOxqZYqR2goXtTuBmahnIDeZMm2yUTbXUEmC2xxG5lsb5QZmxKWrWgL6xTSGtQG0
fs7pqNiuRR0gI6KrbsrjTtyFZqBtEAp2j6BDx10tst/F2dzsG2XsC4W/cYMyNOvY
SiYUzwngegL+AaIUKdN2f8oPeKOcUy5JS1BdHMaubdwHqXi4UCMQ3rgxYo5XROHc
KPjMpSPq7AMx80G2ihNB5YQnbxX1VuMx75IWwAH+vautkuISqyWAenhu9xBWlSol
AUicPNxPqDalEqBJbyT8DNcsP+cAxNAHkYoVGbg7DKPD3hzi/9xRjs0k/CSOBcwp
gfzqW5AeB/8MfGzcW5R/hU8Sg+8vgrcnKvdSiHr8c921kskk1abFRMbsakZM16y1
RxZa8G9+A/fsgWUclTCAhYx1nQGReyrmUQkOeH5ml03hZ3ocIJOWyufG6OvHOF3f
SfolfFT/XyVwRnL0zdXmk8a98u9Ofh6kscNW2xhp0qp6226e3De5uWf0Rz1vikPh
ucW1PMeNiDyaxeQThMFDyu7VTQumbNKf6qzLbr6djvEEiykIsVNhvuIaEZSWJxdr
KxkolIvyAN0ES8WAFE2b2vQRwnbyEoBWBBp0/S21MMVj5Yrz7tOoA+znl3h0+v1y
7LUZ1XmeH+hhCWIYd8BW0LQdS2JduccjmnJ1v7xfwPsEssDnCAx63cTXlK5+KP0m
iiWkr7+B9/wy7HaaA5fW7i+DwfxgbJkaXviRCrO+8ECPzgJrFRqC8FhnLWJdBLL9
0NAZIm7cQt9DqX55g3AwCuiXRjHes5d0asLLMYWYImHRDtY4pnBpCArkiCAdAgMi
cnCAElTV2MryDYN0gLYU15P2+jTIm/CMhzODrE6SeMJZ+XKXaJtDMvS6ETHbOh4u
HElj71azp77cLPyFGkRplbAEpvgrHxlv44Tc/8rAUqeoAWl5QalqzeAoqlAqrVOb
jX0gizhvcqYBI9hZ6sp9eb+OmfkUCT/p29Aya2w/pYAxiGIzJ7Ei1iKJXt6L+Vlk
KBAEETq3o1X68dErIN5nNzbzI04UbRMbKKOpz+WMTA1Z58mmQ185Y4X3XUtaRhHx
n3R9adi27WrNLtpBY2k7+/zuiVahe+8QZ2nmjbilf7vuhvru+BHgHXWsQ9JMBVI+
R064TlN9j8RjKF3jcZlaIEd6Db5ipyhncyifR3p+XiF5aX94YQQ5///bpG7ra2Wy
goWDIaxbDbYR1RKsjxC05K8lF3jG+da7p+Ncr04n7XeHjl6g7jY5+HC0/7oPOmzh
R7tTAWlukHJKlP3AMwKGL9XEzijsqlxx2jdMSUicAddW9qgMCyddKxk4Jb6wRpIQ
aY1NuVSxhwx13PZ+ixt8kgZuFRbNilvoEQD0q/d5gKEh3LxEp2EklJLX70SosRL+
UuUJRNUBwjDaf6YZ44f9EhIFx/0slI98WtJAuwjW9JgDEaNripjXiZibNNA6EVAs
wIMNp013/TWLNnRKazHXr9CuiykB0uffdgNZBC3TsT74umAgMK0+KhpRpQiJIQEB
x2KkMxHWMJeEoouMHEY9y2BggFz8l/cFYb6pZ/nb1qqsTTSktfxjQiOYv7JfBchG
a+HnfC5rNaDVbs2BCaPos6ofBFkuxWd6JXbokOoBvn3jQgoc2pfVFHql3IV+uuED
CWG4GnIkCZ1DqCTnuMtRk5IL+ssXna599lgULJJpjtm7AaMmiwKYaZsIzyQIYnqw
IaMhSAtDmsqwS+sk4UAG7AEGu28uK7ZWgQ23fOklxi5DjEjBqL/aRWKo+p243dCO
QUhZn8rgnINXF14GTlfIU9KbEGVVm7LdN4yLM2qIjo6kQ/BQolXVO7HwNOe8G/Kt
xZAuf7k9yvjd0yyy8JjQlQjk9Z45kKdWoeWjdaGznVjrdAR9dHNzzSFtlrgGFsZz
biFAQnSf737Ts3ksg0PUPrkF77Xcxv3fVOr45RfC32gRXcxzytoZtgNi/3vupCI2
H22upYAWj6L9lhE2lmJKosnQL4K1UZGfk2etUdLwAhRb+axjQTq9Bs3KqGb0uxzN
0moF5Ro/LSbnBtwuDW/sztt6LBUKLrBJKz7+Bch6meBB5Rw78Acq31As/Ie06I5i
wAR+anAiQ6jvjGfkymVM9f1GifaxxKDNMTRJkqrlbmerFgdZAIJvK8iPjLGurtYP
gRWNokjB17sFFRQ5jS3KXzmS5HfiWTUPJX0qGbizgnuD6gSdhi0T14td9C6l/9qD
fsKyR877BOgy3rpQqWPaiSnvqVI9RoZn7cBbHO0jXkKOrwtRFrKOZZF3IJo+T//9
JbWhPoZk13T85rFVK5HCZQ58GVKhm1JEXle+UW/f1IxmQnpyChZXShV42p7DC2Wl
xZtq5Bc741R+H9J8eVLwCMZCAyRoNl1C2dcKQcfzuSFuuLQ3B1H1XExQVKET2y+V
NzDQU8C65E72NIJBHuoaUskK/UlQ8Mmuh/4c6a4v+dA3TQwzC/EuJU9Xi3hylK4K
ZBgEKDXEuK36So9BPQy+Sq2APiYMi2sMPBl5wmnOHj+ZnOyZe30HDP9NqmS//E3g
hjA+g4CjkTCP0iBckdB5sWobWXMr7KXss8aJfTJbmClCXW/YdEgV2f5oiUkFy5pI
a6+7bMhG2igvAsmpioehPreNt4eITo27TCFdr2i0dWWkUkJOP1wugCLazhY2BNnC
r1hhKzrk+hCn+1CuT1gmq+l0r1mYEuEBlvIKWrRtaQVagxkgl3VBPqIvIIeQK32v
1P9kmYamMmVJvb1mhfxIHQMq/HaYnUpaUvrUtGEgP6UJAfmCJxUHBe2eEr09R+vm
0qH9jNMTj4K/4FcX4NYlT8h4MSRW19+iXxCEKJj4nTamgL8QREZPJ5e2V75AZvcZ
xP+S+fwi6w7qdZ/WanJXlfBcww0bZM0QyiJlOXkR3euH/cSrvBPSpEXL8jxS2Uuf
TaSUrRZ0jkMLZGtNEdX8jKMXGWM8zq+FtqKu5Hg9lCU/WdlMJzd9XnC5URl+gI4E
77P1syHRTKwHh1Tas0dmnHGfQeBulisZzVC/WxLMU1EplaHkU8kFl0OE6j2Y139N
Lc678Ftoju3hszMlwyjatKuOl6048tHUG1NqRqJHQnTjHdXKHYtQBsiIAKJEMYbm
2HviqfhLYz8mesMlfCEFqJOTTMoAPmKOXwL1VrxmzaW3N4JpCpuioef8RiguoIzM
82ojwYixBECKM+p8Gyg7yuNgZ36jYln7PASHf5OAhBv/9o9saYoBVHLtcEWZEfsG
7iLkI6kpVXhKvF1kfxdKLHmFIYKvEaY+3L1HkLZ9vIgRodO8kaMAPabGYjPYOSZe
QokdzRN9YrJ5PtqVy9kV6F2uR95IffcTDa0m8uYBFPJZqT54YSo3ZltqM3WkvEe8
DQjJMzaq76cfZvLUCFrPZXTTgauWTSyGK03/zY/3jz0Prj6afyxjZqxOetlK3IxB
jBFNKS+e+FOS4gg28qAq4XAOnS0l6YjW/Z2DKaWMF7C1xb+dpfrAVwaeWaPQdXfm
sCWYONFkAZ0/FejGpNnsI41Ccfp3OD72R30WGoNLJmmAs3zIcgT8r5SJJ6Gg49Nk
SNLeyBtVSF5Q5NoFUvPjoA3kpjQF6MFhDeDXaIwbTZYtIjWKv7IIpiS04DyQVgpQ
vl1QG+Bx8Lg/BDyOlCzVuzKXGvOEyORIY8yQ15nIWFw9D1r8BCGlE6i6YYK7WDqP
+QgOe3k8UBpP2sNJ0p3AOeAyngE06i5MP94a2fxEW6vo6mmgQe8uWQq8DiDcG+9M
Hzy2DYOwcfVJQzZSJRmyET18PZSwt4nfcuvLjDBKfe81SnLoQPq+W0RbHQOQEJFQ
UQIbhLZhb/cvhsKbSLSBgXf/k1zzJsFrHO1iTeb/BWBmiQNPusrTo4w/ry2pDAsw
KjknTwTn/ae1z39kNE+3An60bYRv2WHKKungnen6NpDzwormkewAUPPdx/1x98Ja
iLnnkCOcQ1GvNvSJ5pQM8iaUT9bn9BEDs4T+XvjecSzwl7pmm3/kUvMF6ZvZ/jBa
URkkctXVqgLegOD1ABT4WKwUPn9IAap8Kb7p67SEuTFBIteKbXLpnlcGRfgsMUU9
dTIDymm6OFaRD1GEhH49u+6OjStEYHkCm4Jz8e3+d2I2EBfNBaVcxNfqwWWfFfSA
oIqawcTW85YopX21NBdzsqHIrEZQmgsmWgkunLq0qR16/En3J90Vixl7dd0dw+z3
1g5gP2I5dIC8WHwkpVAxXyCLCKYwLtFHHFAeLlTmqGJwopo4hIkVdJxz6l0Hl3V/
HC/6Xx3jQPIfcUSvLGZ+dr42UXDXvIVHPe17iCT/BlYsTaG5HlOF8AQx04VB6OPy
iqPvKCTvKiLZg5nfTG1NSdcJdBwVpgO9LFuHMXuNLJa9ZIVf+DNqXqONvQ1TIFjC
OkunpxVrKCqJPyCG+uhnkLRUVVI4vUBJ0VcAieXoOSQDkIngXjTavbWW87ufFBY6
AyzGkGqKq9sgE0X6Hdj/aQXEQAaKNrvtRV05PAnG0GLX+1M5AoH5QW0Pc30N7cVw
BhJn+c06qatzotIy0qHA7BlEgRymQHtwUkF7junZrmGyplXKLyyov0QQwIJlM2jE
Jwiam0TuH2eHXQJ22Vew0ZG1JVMNzqZnu9nNgE9Bv8/TIQ+Dh6MBf/Iua2/ppkuT
mA8Wc5QaMmKernnvw7l3WIW0uQYZ6HB/K0lM//rz+T6TXGNiQ9BFbOcxoJPE47tO
l/4bg1oxpgG+lTzLGMO/4nyMzjWykj6UAhX8nbPw3/dSS17RugO9Ps5rwJUYP5xz
tOE/MaFqtd60qD6HZe+y0E1P9744llz6tyVKQv8qem1wXkzITfmbDgJN0Y6z9bt6
agK3ITmwaUTn2bVg8/n76xLyPb1c2YQXX+zZQktmyEpm8VN2UcMup6oJxxFND9cV
p4+do+xf7NzD7stwdlfPKC3jdy5cUUPD1GMftyQ2MYtHBc9BJrhabevssCiUbetu
wdlb6jZNlUnoj8PtmXlYk70HZkY+6sdrPNJ5y5YcsDHHlJaqAugTn5MDqx7W7dK2
WjM86B8wXORPgnm3dEwt4f3O3HX0Q4RTmV0uCT4CFHqnCYweq4TfMxaip5tfVIRw
y3O36BaWVeoeUYrZYcEVVoEMW0gL3E9McvqyVmZl07sS6FaDyRgC3B5lmA+Q855x
CRje7Skw6KbLJQKjDk6NSR5tPlkWYHAblM/RFrxONmhUwUo65AMd1DrcO0WFV/F4
fpepJ6yjZ6itR7BxStvlC7BGsXAozX6sKF62kUHEv+hVZeeW2CEcjoQXDiaxv7bs
81+kuOKuhAnwrIeMDMT1fkEQ8e/AbzAew+39Dccr+EvF6iY37steayoIxSEQtdrr
VSuL/Z+Pyys6w85JWBPsdJd/KQudp5ik+dvR93tZzUJBnramebPYGTiv4/nVeF13
KTsET7n05nYf2b2cHQVeXHzt7tkpcTflkSRZhKjkF5nheiq6355sqTWsxWKUejlC
LLHtz4NPH7EieeTbpqJBdGFE9nxlyAIkeyl/KbYDgLDwro3+XoXo21PsDlRkWyAM
WiZp0NHb0PxCRRqIBck/TEfgjkbTmeD5o1HvMl7vephwx0YC9rJhNx4YL9DYPvKf
BJqUGPdDaA7hY7pB1blKrhQZs3yFQNYB/4s7N/lhxKCKTzfenoEJs4IMhj9h2RI2
O6TZndhJVn+sMe4kCyDmjJnfCfyVl3E4ziBtyjQMNzLSW/QkWIM2y8oQcRuJosmT
RAGA9mqSSc+Zvi/puMb18kR1JBhKOjfqIzhKnzVTV779agrVwshHESGwGYQN+/7u
q3A19SVJD2JC+6lYNBXwxSVLt4n1MQIQkIH3DCWlyG37HGArSoYnOvIEKKny+ZsM
XyZboLkoaZz46wsxU8MnIUlrWPCo1jVdNsisvd4SVUech0zEJbh1I9qe5/6o/xI5
Vg0Ypcj2cTipReYIPjwYA+L/J5bl6i31Mnpv9QHtj+wve88YvByOU+z/unTXnhFR
o9gUFnVaK5EKw+Mj7IzC+TDzAz/G/TpDFo37n1ObwnDHcD/kBqIW2urcLlVUn7r7
svqDs79fTHfLo84f4Gw7sKMlplhGPxA4cI8p3xWL4sP/mypUEV+mXfNdtTSwyl/Q
q3D01zlGTxeGKKq62vd/QEzLwT4CMu1MbROoCHoFHrtwgUBMMl5sfwkHeCuLgoEz
4EJsp5mtncG3uUQ3PI3gQxnbN/eyjUnoUYyCNpk3l6+DzNV4ZJcaaLtT894tiLa6
c/l9AeIiJM9jAdQeaWIvMMVG8NHG+3EVX/b67uaqqmisqTy+3ZTCgmm5TEQO3YSn
eWXoK5TD/2ZBXO8V9UunYQUr/aRtSQf4XkOd0QuTArm7B5s60bO9Zjk6J4x3D8Wd
sTCR01fCASb7hH1tib2v15nq/0vrPb0xaWXWthRxqoS/0u33EV9iVt5i0N8G+r2A
WT9jPwLqwYQcjc+Uht1tJDQHa0ntmxldw1l/yg8cSx4EfDfLN++lyv6BMoHz91AY
lyJ+sUEENEpaUT6ZuIghs1LkPkL8/7T+6yPRja+moBiE8pqeqlFHiy7QwbpQplUr
ArlVX+B1FKhemAoKGWtBD3+cHv243eF5Bj7o8wKmXrpvF1C9BSO8i7+KqNj9k2PA
32lo4ZDpUw/pg3sV+xPnMZeCnG6U254I+PzBcCmQAxVG4/EzOm3WQbfbmTtTI9Ru
MniHSH21M2FEL9fgKHp2J71Xz8wdkpFHoVQ5MsIngFXhC/T6XBgRdqDFmMTy/gzp
KMtAKK76q3IhGuB4NxXwxfpdsy7V3t2NietkqY8RyIniCtYPapyw3n6dOmt8GmQD
CaWuqImXMACQiWas5gU3B9bZ/VEJG0vExRoFZukNX4UIr3eMyQvtzVJyqzDZTVkZ
hKkHu9cf+8JFaK0shEKXIR8+k3kCXwRG7Y2KnjGZxuSp56Tb/933oBe4b3V1D70J
BG93qjHkmDNn6eujJf5JeLHpL7kzIFAg6v9X5Pl02hufxlxDvz5ZHkoguUjHFDML
iRwfWlWJ6iLPQxYjRRHqE5ZV6hxvbOa/gh6Swjp6JvEf/fzX1QdEc/Kx8P0i861K
zA0Dg/Kebc3ooNZsDo0xR3Sm86Ze8jgNwRpcO9vnAxZmNUIu75YhYHe9qYd3211c
eygLzsnRWwWgeEq+P4bpTCNQjBBmv3LRfMKaisSeY6Y/i6Skz/9kKR3OpxP3eEok
Mv5BGnVZVV22smpz5tpiGQ3ckY2FyU/D+jcgZ/S99/DEQIWIRhmiLvb07Qqi4ZK0
veP2rteQHkYAYk3jCGgi5Mp/8kzNa8biI8kIKwN1seyzoSerdKGIXIymJoa0CJNP
buXuLs+pJIc6UgZiGIWXRkvjsvm7MvLLpoLbcLpG/RGiETS9OEVt2tgRMYniyQF/
CjrHBsm7tQHnMQJWvsbrhoeqqfZslfhRoDVZlIzEf4ommcj5gpHD8RjDBan4yc5x
KrKSQtffWgRHy7nGq1Xs861RKu7moWMs0wzP+Dh7EW0WE8A5YmjqWkzdpNZ7VqTy
KtNOv0jqizTog4SpctBRiFGMJTeqTRbAt5KYnUAgkn89oyyYVvnaG8XJtwQNBmE0
qQ7KwAWc8VGFHHzuVo433iQUt3OvakuMfG/h1eoXHuzzFsF9AIk/l2PxX9zDWvXH
ah2XXH7so71NtkFVimgaRtFE2pNqv/5GWWIDTpswe0crX7o48EYDgTqRMfYHLolu
1rJTP3/HgbQc0WXPj6TuqzbY7ZpMsAIWTn6fkmPV8EBSsX6f+h2U3B+4+xCCUxki
90UglAJ/AKGAKi2Lhdysyk+hW9ytvFGuYwMUC3C82p+rcG8XwBbkDS24NBpAPdo8
r6SMFC7LeOmjZGSX8EP04NCD9YA7Gjt4mOgALFpOZY8/LLTJi9WIzN3WMsg+ZXL/
DibODwNG0KM/GF2SbItWzBwD15n7VrYg59YBk8NGGaeZAPpNo8mLFbb4fJpAlfnK
cXMQOQqidV+QYzHb2wC6lPWyycucuhCZmb8gx1J6EV+xs3+osIsTI9456JSY9H8w
EjOlVBJVSY2h6RuYgXWUGsOgQ37glbx5BrQ8jPU6wD1Jd8Pkn+huSMfaydsjR9bo
PWqKt2V9g9nLKhZmx1EuA4XsQlVRBAqjzdpC6Tn29ugmkKaZCi6kvlRP70XEQhp8
X1FTW8yoRN3nnBZ+cy2tYI0Y+tdC5f0/jAt2h72AAp1QJg5rs8kRKLYltct81UkL
dVtVO+fMJkFtygfcFP8QGbITQynTCu1t5SgBATvtNAk7vf9yh+UiIdtH0x8YhI2W
MXedt8U/JQIELBQ3TLEC+7K28lrgiiQ0hfW5kW6SCWVEcD8FOz9qwu7QJ87Bw25O
UsjQCVfE0AQvZjevHENXUb8f5KrSANNybK8uI5U3N4vrDIQIs/RtnFsyrkNve5n6
I7jw9X7ytClQPUZEelMA2KXq7QYPsXaj7UqVTAMoh9bZp2+kGJperQZ2uzGASXJx
NU8uWR1qed/DF41F1cJsI6sqmyWnNaacK+8gaaAccsfgiqIEbpCgSdfagVUr1/ga
eh/GB/Jp5HthX8hEsAu+2dj6TJGamJEw7/ZJToGDN66yKAK/gK8nkqXInGffjwRx
NaIPnHy74ErELI29U3R+kiJ/YfG1lcaiX5vsOmNYHxtwvCaz+OFDCxjBysjkevmj
lMxp9Ec+PV4GQmbBNPHi0Qjb3nLoc/XcaxE0e3Kr5OrFvKx/pxPNOdAfBIbW0VhD
fB4YERok48wpEeak5muZTIZuoUCO7dczO3Q761COjitgdyKycOePQ/ZU6L0TiHKz
L5RD8S4rhRcm8zqZ+ZvppcaqNas8gS/S8U7RD88gqKcWsI56BkDM1iSb4eeLOJOs
FfcF1UH49f+6KNy1iM0lAdlRJoK9Wb8ViHXgddD/e1qrswJwsqNLmJCmp2i6P22G
Mk5s9vnkhUw0NWInyxS3MrbQx/3GD3hr/lKTLmnitsFIMdbCSkG2PV2IzDUkQbmi
syAZMaVARReKZLV4L4X1dzDY5MEMNY/N2lPbi15sl2wBt9jeoKBsCwxvKcAVbr2q
YqE04I19bHxV6GvUIlilBWaEUTBt6pzqGVB+jIX/EiQbXU4VvSGR/EitPZSS/Q61
76mRAjkVzRKrgB4b3L+hPFuDIEaAsFLGM6wKMtsl52hgbZT17yUYEGvzd0/N56Ck
XWqkY+tKhh8qdant6m81YTyTmrSlm9EttlqdPA1ExOYU41p1RGKzcG7f6eAFE/QN
FG8JN1rFjCSCJUX9qENnkc9hhZV9HusOUuGMA6R9KWbbBLll27X3b3qmG+YsRffR
rOVjnBe+luhwB6UH/jKdAh4OpxYHdPPY8FzjbAlD4PDe0V2ryfGWlKjBThMes6us
f7AQWXV6lJ22Ec1RK8Lr2P06XiQqLiB2QrCN/n91KNwIIlAkJbHWroF1HyGyDCdj
UCiLlT/LeGD2av3KGe/bbvkiL11kKnIRFEhcUF/VBenBO5qXHTTkrwoteQiHL9Th
itccrPilTt5nl4aSlLPWk2PmJ/G/+GKjx98aQk+FnsegOW763L7hI8RwR5luK4pS
cmPozHCWOgatp1AmPuPmSwcIpV3eP/q658YDTeZRYyaTnpteXQ/b55Wk7yzPXxF8
W/YKqfy3bOsxTZXkFJJ9gbxAnsIPuOiM/F96fUPQU/ukgoMZJO0z4qoMIz73JV11
mszzDYZJeDaKxpdNW99zY7u23wz5pEz/NSgnAN/53GmXSuijaiM+Bt96sIoHntXo
OD/0V6SiWBv7l2XcPFjCnUK31ratBxJtTJjsDyo4l+GJOCiG/s03Eeb4ovImwW9d
5g8t2dxTZn92B3jNzWQ2YcLzk9O6UqyaaJMwJZl+GD/FyKzKCRyL9oAoxPGP3ihf
cs8ahnEz28+xGWbx0wwASv8ey0fB5MWNeVeW6aT8B1Awm/NNbRS0/evt43KiaiFa
+Eyyszdplt/Vx/jYpnRUf8GqpYYq7GWi45UdJgS8lCqN4AI5dkDzAROpR9fchhKS
o1207j6YjhRnmBqMG0WldNKL4RBT0k+j6P/qdoxe81C9UsGqDwRjukBXF/PLcCBB
HXfiR9x+IS5OPMSUKGrNUJ0/KfIZ7EUP2QycwOdfM5iXfEp0ALbaROd+wzXKAyFV
XnPSjqvGfjXufZOp9Pfewa3lLSJlflcRL1ayPnGIlj+HvzOZ45JEjFB62tP4hQbJ
IqOHPIXoVKDo3DwZKB3ZiCHBVpFw0v1J3OcLH4MRJVww3tOjFPlMW02Ws0SwX2/v
HXOoA5ql0UoQBizk323/ajK3adJgjt38SVoZOjYLdF8a+or/u5mtU1/o5aMjXeKX
F5jTbmJYElWEGE4l58N+7rZ+HnK3SiONTO6NNHFieUpCJxULYhmco6puvVXrsF+U
IpLTuyF0kndjbAYxl8g82MVE/S65+Ff56epNFuKZpw38AYMrCNnEbapU1NDM0/G8
BK1AH9/S2odISZ/cW7b1s24xfxT4Di8/KX6kelulFedLIYJoJOvfJQpb5atmLDCM
KP9KuIGpJivJKprlgZYMInMvB3aRuGt87Mf2QD7Lht7a/uZntNB0HwLKNGuQKhm4
gP9GCeMkMDvYihLAgWGRMjrqFgY/XNa9RoxMjRivQ+61pTrW2knMl8Qcsss2iSUO
qHq7cfOrHnq7bgxZW3zWihQYcD0QHl1FZ277Sb+X2l04daaxY+iDQb8ypumflkTh
auOQzV/kz/kqCwuk8mP2U85arHDfse8L25CaII9iJCDoxcKaKElmXKTBH42bmG+4
ruvZ+oVm2KMImv6aX41Kz81j+a9rBl6UiuJg8c2xpqG3g7tteJPsikAelm7fepNJ
mt2RL2XruY61oXMeQFW6o5RmVbsJresbNra5oQzU2dRj5tl2pfW2km2nOTz+c7Ob
wKGB0GDGgNL7Wvd0IgCPn5j23ASGefu8A+jJ3hb4873QV4MDq0+qGQ4A2/MAWfYd
WIdAX24DYxiPl9KnpbUxo56sYAwEEHJ+i9bjekgr9CxSvTvItjwxthKt45rh7Glz
szE2LkTUzJIFdoFD0tGcWwQ/9AedUe24W22TMpErILhq9CNZaDCz/e8UX0sg4VdB
6bIBvPMsTG53dWMe+87Z5cMB1R5GhMtOnwiPXMD6CCuLJMZEytflzvLZn5FbQbp/
KiUcTUvlZrr779jWElkYpR0IZOtx6tUALZX55sNJbFKwcfG5BEPp+O3dVcdrZXWZ
Whkv4566gXW0Y3yU5Bwu5kWksUVlCjQeTXKyUbiC2wKtW2Vjo2H9J4n2kFwCWDXq
tvZBYHwDZqHKchQ6sndFfP0EC20APsiajzKLvKTb0ccoADnSDs8f0y6/nZgmCwB0
uPU2zcZfkSSVt3gfH9+d5TYDg4gPsNCUbtO2cVrdiL3HRkrNNnY/BZ3Tf6XU9hGC
yyAdvn6pGyVLAvPgzS5Wmk2kxseQvsx6iECLieclLeR80qJriOVhTEjuDHBd5yON
/m+3liCejzUrnwn+IrxS1/bufgnFLQfCIR82YFyOJv16dTwKVNe73XHCh97caD6N
8arbm8OSkpisyF2PJbWWlee7dE9yi2F+fxPpTvRdr7ev2H+vb9QVqOKYf6OOFdXz
zptvjcgkRYULqld3JEq2H3h1N+rpmbzfCm+Ipk2+oy9bRh3qgAGpHTwhNImuJjkI
5DABgZpqp7G8+6Zq1DWaBvQESAMVpkNYATKQFKYomXFrCpvs9VGqEQizgW9nFZIB
xdEH7PAAcnFkO7Bsj2jBA2qXDvciX13/fSn4qLUOA/ixYyg0Nm2+sbRjhH7qDSPe
Zm3ZOsp3IJ02eaAbSvtYRyeXFx0uPtphw0cV06jDmIemdWLUqOrzos8VtbIkbxGr
Vu5VG6O+KEhhsOWH1PSl6GfSh0iUJ4c020Wt5BOUxh35jFA18FqGWOpE5jWYuMwr
`pragma protect end_protected
