// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:39 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bKaDXzbslt5Oj5S2QaizXw8TS38KBwRZXcpGnEyHWYy1oAqlmmaYm3b6m6FHhEbJ
qyCe0RPgrUyvbcjU2B9VqX5aVv2p4FeEqlnrceAHgLBRAMa+0Uq9uPCkqmj51svE
yM2xkOcg1AYJELhcTPn6BVReXmibNB7/Z6hso/S85ic=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3792)
akN+nxUyxuEItxFxlvZdkRhvi2Ug2+EhwqCzgvOjZIr+ao1dRsp4e4PgRnapvW3M
930meUyKXParWJV9OxcVSgcgdGoZMhDcHBdBBejI3yp4/3lpSKwYCnt6jcLi2UPh
++ASJp0QBdVjMIWaPcXBZnY/2RVXwf39t/tgf6MNaIlIrE27DgpmOuhh3vbG3Jix
Dk3isDo5oqtSuWlc0ZSSFFX1Ii6Dd4xBujjnu9gshR0m/DwCabwrQBQyBxz0W6c+
FXW6C7S0GVhW8EY/txVKDqPb1LvTLrgT4UmE9Y9hPeAFYfLYKKaVzX4TSl5NIQmN
+L+RMzYm/+PWGNKpBLoRZAc7GWGZ0T8ypJvXBhA1gUkqu6N7j6dPi23OfL3gUhcz
adbxxYJOxbUKLvPDR9CulD13a+RzpIPKKvmqvRcbxSTjnQ+8CQmnnUi8rfXLHSGo
23K4OkoGG5L9aniF2L/wbwQdtklSHmuuds5IqKCiIl8fQrb2au2F4ADOGWncUjvP
Yd0cpYBGGjuTUJKMv136kpPQUSoWcMFD6GIzRILNM28OOdKJI3WDZT6eYSIYERZV
bOxyVok/LNYEEZK8YtMrp9EJLuQAWCEn+zUNy0QJmrNoBN+HCe1WUfemKzqujn0F
iNMaSqi2+D6LiUVl6XPiH9IWDZx1O6OzBaCLq2mexP79YQ8Tc/TsD8Xke0kyNmtM
7KMRRd/gzS78TOQbMnFIjwYU6NBuVkOF3V/On2Fbdl8rZFN6PUMKyYa21zy/uGQ1
Iv+rCGio6JWMeSutqVaX5P6RZ8g01YtZ7pSOgFGEsiq2CrYe1yJIHkDzZBUT6QqI
yhwACWyOb2EnquELJIUpv8SPDCqh9m3onWOZVzUuW+WG0XwViKmZs8gjxL4jHXee
8lyMHyFRrBBnC6g/gSvnHe/LXnRkfZtqFhr0JQvuW6ggLMu50qAYgan5OrfUej8o
0LjccmPDL90WpKyKjMPMmtkG5C36u+gOmgHskjppzXJHt/o2diNjbenFhQ4JLlmM
3SIuKTcs6HAfve/te+TXhCSXyDGfN3dDG4+yB9YLanicOm7UeDIbkVSK6tUKTey4
deYEg91Q9mBw6JUQsUnhIFfUQOnI+WJXukS8XoS/LSBZGqs30h5cJqNJMsWjVoum
RRsOMb17lllFSmqxjQjgV4ocr5a4KZPFht9AlrV0l1lKAIN2IzO+zRU7ZPxps+Pg
3j6KE7npU2IVDcjB68cIhpiheUVK6wscTocNdEBoS7dip+wxAKrxmcQOJNQEPby2
8PKx6PfHp9in7VpEjSkZCkaw8PrvQ4sijfMhwilg+jUHQsuiroGmxKO4z4qzIr26
pgoM709JP5lIGZTmmKZob3Kf10jOzQNlv0I3bBgWteSGM24DkVzzkrC/h9iM17PQ
JVmuVH7lrArr7LGb4olWNO4Y4pAaS5hwdsC53Ciw9arY5r+JC8VStL58Ts8CqiB0
lWg2GTZY80ht/L6AYxtNQ2+N7SOY1wfbFfcw5csqKQN7jl4bytg2au3H9apRCR3a
62QOw38YWbRAt2VGtECZNadATjqqJFKLS0YVKbCyTOBlksPziydA9wrh571diMOW
dm/ZlIvwiCQvgsfhNwF5TwaVL/WvCkjztZVhfXGAuoKDTPp5Q5zyyVuZjc1TJzZB
+9FLvzrECuJ1y9IodCoD4Ugvm2YtpdJJuBg/3Ksgdj0keoMNS2rw9W3dM34Spz8i
t8DowLbi5f1dpY58GL8bDkJCCw7eYDFB5nIbJg2i7hP8oJxnvVkhJHEGkoP3f85I
CeIVjUrEkddHs31fkB0P+wX92hN2OC+YEjO3t7DcqJAgdnyAEmn2+d34CXdkvbdN
LEYd95HzsaZNvFqVSXWKqlmnrH3B+/jkUf4LghBQ7XlcwaWrIxaGotZvAdfCF2JW
gpX2kiVLznbDmMk0FOazt3WYPW3KiEx53HnOTff4Mi3p12RLXkJqTj0Qdccu+i/z
MMY2D1v4dIX9/uaLgMgsgEADnE9iX+Qor8Dkqea43D9/2qjPcWDRviqTxFBXw4UE
hb7x5oFvUnBprpIiMeOiowTYd9ihbMwgOH9K9h7FkGLDH5cbKtFVs9pM0zXx6pq7
fMpx6twk4q3MFV1vXSGHvqwUxSKy0D6ZjWisJ9QPHpJ9AIYMq3OUQ2a5/4e+kWaw
O1VE1m6LpIK7jF/EnYREkDK2tuOv/m3Us/YlMioPmiPCIvGi5RpFvLd426LaO4zI
wIh/8vYcEMaW7RQh/0Vi7fXZEA37pjORD/4i837IDfOCNuL6Rs2ek97lmRr/Tisv
wM4qCPty5SRB52g8SVO1Bh1rP6SsvJaZpu/gDW+NdVTq49nUI59UOUpSqJ36rCEk
AFO76lwfvb5oxaQSR7SYeE6PgiBF/TmH3M9cg8ADDWCkZXegEQuSL38NY3GZ4lMs
jq0cmcf6AzgBCIP1YyQImU+sXEFrZUqqtk9t1Y9HxQ7J4vuUPEKL3Wae0nQAc2+X
iGgwg0CMVc9Ap+hMuMbagmBL36xDqEAacsip7I17JAwzbUzh9UC/jhRgK7BDjyRY
E9oobOOuOFopbMvIrJwK0kvVCKOFRws7Pors6TrOkf4sz6ckEViRu+PlXBRiD94N
8o2eCfkuKr55DtR5GIz6+l+BTaO9LHPzePdnskTAIbYhhzu7YBjf9bpA5F8cbN/B
fIN/34NbV3P638MP2nyC+rlVHprdlJSFoulGH0JYQtvxu5BgfUxpOuRdPBfy3Brj
fwaIja1sS0WpSXehkHP9XQONZ9nncVUbCsvOvNL9KLgKyYzYs9TpXLS1whswdZlO
gejDgXqp3kmLndKhQ6VBo+iVJ8aeo+YY4URbFZ6UKirdb+rAI7Ki2TCJQv7wTdgu
tFE1c4dr9UnQLmil9bJBbudUSGP4qGSQkZLnlX1II2599lRr2d4ej3lGpFUelaGi
IIw35xbYm52imyXCZFraOlKfCRc0Vc/ss7KdJaPlYO9l8IlaaN25E116jxLSKVMH
Wmp13SUXp3GoT1/kiccmhr7oF6cH2PEVWU0ZClaR9kCmMDh2C8ys/+IctEqV9/dJ
F78G6v2vR1kbb4bmYntrOgMq15zSLodCtpRV4WEhDfIZ1SDysbjcpzHNC8amrqd9
cthcFUoMgcxBXoyB4ssSs+JIQXr8kgxcqtQoqrwDrh1iTRWT44/H0js6i0MSHeWu
58pGZOk3UTvDqn5CW1JLG7nYwW2Omso8NQ46R7yik+XV07ONMVGYDfcKssO7t9l9
dSoKPca3mS3OrD32OY9sYx7uXHrvfYE5lBqru5bkfJ6qunKKKjujIZ6MXJlQY2Dh
qrtFxD9JMaX+cysIPt1Jr6notErcL3ggaLooYgIAmhhwlk/6B5isuM+vy1573wML
V01v2Iji5l4eBJOtL3iBA2r31qeCqlsb8AYABIlzHO5SvGTnPXwkelWkoxvbaArj
V5P7xlNo178VIuymGorr5Yv9HUNhOqAuzFfIFg0dVdrD2H9w2kdBrqwCgNFi3iLN
8FLVe2Am5/saSp5scvXweBD/Edt4D38cFExeCpNWXNPvl65Ymp3BnprDsspImyae
JPwdJ08FNScKcVOqL7rqNNfmvJ8uCLa43YevIgqlrQyyi9KpWFQgCeV/Gg6nYdSd
zKsXc/8BDg+WSVfSPD096LZ0g3Pkz2utn46m9QDe11atf8N3Dg0bHwy1ljpIhJTR
UXLuJVwXx/NOStyM3FZK+o6biMbGNDart7AOvX/W8yLmxxYwFQJBTnQDGilwJ0/6
Gm2MZPp4d0Kte6eMyteR9k1EBmryOe9gx+dObDeW8WE/SKUo7T0P0HMNqoZjSc1J
woeehN4FArHJb5EerfMDYWVeLYtZtImpAIcPpNOLRunoNdkoqMBNejLdMFTkb0sJ
/oHZ89lQxUB0EBTSF2hRR0a10Vm3Ygu6wP+eF/UMb5VTU+/olZlZoE21tEIHu1NV
qFIHpEIP9mYrvsLn07bgWDM9i93MkQ4QTytAZZ905rPhGEVlUdSyyOZrrtT7YZDE
dUvQ+3mO/6M5eWlMymq9hHZ+jb8l+H7MGMSNmDOy+wlyvGexJbYTJAzP2i3lDwVr
61OLCRbx9dEl9AB4Ljl5aXorTEHwglduK0MkvJGdwT6SW72CFOSGsKIF4lz4yPFY
km2qoizzPuTGo3RpKBy7IzBzIdSwlNkiS0p7C+UWMAs/XKj4ZOSJkzn8mIDXMvSC
PQJ6WBkkNJUOcap/fgc1bcrOe+aGVcsieDkoKn3B8vwWhLEh7KKrKWUX64RmBh9Z
C96mklUI/X3kO7klwdAXyBniYD6whHQsVwxxoQylDCTXbPet0gbAYWyz6xzD+dkH
FURmWxSzTBcNcVgA5iscq87LIvIyPbNytRBqWO2e1E8nhmL7aoqvGuh2j7LYGRGu
BkUNuFB4jh24aleX0yEquX8PpSlL/10BUaBzKlVqI1Wh7BsaDzwortc/umCDDkON
wSyU6TsLuEYLVKMej5eb/Jyt4sBZX47J+kX7ljSyczTVeWjHdPTP0jWOkgcfqrBI
naS5of+W3Ap33ZpN+aksXifTnH0OEDsTqsyPxfDQWZP+wRv61oR+wSg3ptdC7hmS
504fFTl+mT9G99m5gQ2KCXeWmIsg3PpdHGnQOeHhzCVD+FHrFZX3GJrhuzR2jxAa
+77nMWvGghYymPysZxNaLdEziEGb5LVSxuAqyWHu3ZT6F0y7KmGauQ2d3VnovDTD
oipIuUdOP1e3CA3LIg9QaknGoweovObiVtoR/ZFh3Z264BnJmRRNv+SQMmHOzdsD
EAsjo6ELv6sTPcZsQ0zaKw2M9bOw7MRpxoYE1drD8gWd/nejmegMbtESuav4Zofn
P1UkfYp9D7JNRJjj1YNPQ16j8krcf8bDQI24xRt4+yDGF3zNRO7W0J8dgYffSLDD
b0IJj+nWN5hh0p0R7VaMTLXmJ82PBMYPywczAcy00hgXCf7PPfE6B6ol7oHRA4o2
5nE4/Rj4QsOGjiPDRTj3PxOsqCFQWNO5vXCcU9AAJ3RMe/05uh6YP9cn05/VVHgf
`pragma protect end_protected
