// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:36 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
T9KnWaQHBhCJ5kX2poZ0gHq/fBLMYyFXJLhlSkPlXB0KJdEziCEKlOtZDegnJfAT
UI6bdsr853vZnGNa5B0BA4ukLRkIXEBRYTCGpFbDLhSpaTwc7vyGZwOv3+OBWzQ8
XEv//AdTrcFISmu2Qu6FTwXdATK0WpAv2gCxp0l7KnU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22080)
6ktvMVs7jDl2KNeMc60wIIrNPqNgubDyWeUitUeSeUyIwctNFMOlc8bpcG8UBUyl
3lNFyNetSSbZrLkt1qpD5yGqOWjMUj5l4Xjy+MUeXwJVNktcDQRFBGtJWlsocknp
MhcHHuWLFBjwqpLK3tpfcOauZ2PjUDV39jfdE13kMBXdTIu5RhGQRLwLCHAm792V
9PINjfsGV2I4PghCxz7p3loWs1HwiK5SvMJ0he768o7cRxmOBAmfLzhxlBJx7abo
VfWA7VT8U24nJ719hloxvq9GMTSRzIGMjchUIY/jc8L+sjYLAtg24fe/s8ynj3Fi
LR1Pxyf3M4ASk4RMkBGz0r2+/RCY0/KowvR9me2rH488gdY3aV3MuyyO2o/A/0R6
xE8E8c0D1SLB/SDXX2wzLNsOKyCu9Io/EkKEg0cDd2wPhkwSAUWmBlHAf5WAsuuG
IVlKxskH/aVsrwGDB8+cjC9aJ/KB4JE7EFiyeiFoLmPlALh8ivTTN8lzqNDvYJK3
5Mfq8R8OjQQTgTiAkodvJ11EEqiAcJ65DltXIUS05SmYU74Wy0G9iS5GzFqtuQCY
hUYlUBaoT66xM/qmpCuN1/MansZ+DaILs9hXZZ7/EJg50IRA/4nlEJvohpYBHIs5
rQKII3D45yrR8lVAsgtOyBztbWovBeQO3Zf/VZc3ayiCU+w0ZKMJsu1Ac1L4uyRY
oYZNCmd049LWdr+KCPdaxtzlp/4LJEgaoypY8DlwC1stlm4rOdm+nlop55+HHg6R
VYyZDJv2BlflZvkMQBALF07Q8bhDO+CzF560J9sBNsn56FwVg125NzSaKVrYDrAu
Mujw/EsltLz3KrrUJeUQt6grGRdXYr0tsI2zQYP7rVC9CAUXzBn+SZNIjo48gkw4
YpfWMRgLhsON7RHXngzM6xsBtriRa7BKnZFwWBW41VhtKopZCbrbj1tKeqfuEkcO
GKTX4JYY7SQ7rLZ0Iu1r9CKwVdqeVW3qd8kdXn7e/JlghyNhddqilxoecHP3IQfg
tOT5OdqsrgFJZbpa3VNJKHcItVb4fueTxaIHUUwQxzEJrCgWSFj8kX/EoJvW3zvJ
lcY5sqKSL4ltloLpAvcJTP+7TP0JI3gy1ipVXkt/KeJB7U1xNXleBvarePmOJTS4
18r2QcEA1gl0q0XvM2C9CXYoJJJJ16aI+FSxsynTM64HEevHAJrpne1Z+xOSbdwk
TjAPNIf7X7t2eMZFSgnXHNmsZUdt+KdpjySMZfoLLgSZcwnmnjyTuH5CVUopMDbx
fuNWtAvxLd13dCwC98DwR7De0WR4w8XxCqZBrYDA5gNh7pFCIvIcoQiDtgGBdugR
Gr+OvgVMOhI1vbuiHxgFb0KuuT9AewCGipcBiDKoyKZKtMB+j43QqC10mnEhhDG7
lTr7DFZ8N4wzY6qJkyPDBZ3U1XJeFkD1vG0O3Gg5c/2LOOz3HVSFdCWIwNdCskIS
os2DH92RtEQ4imTrLxmfcS/ZuSGDN60G7+ZxnJBUdFWjGCPfEoxxEu1Lm/UVmg0S
TwSf2NboztfdDUR8ezxEL7RqxKbD7OUA8VdlHEg/y5ZkpW5eHV+eBonWRbPL2vGX
+dVO+CqTitvFakjT9f2qmq5O4FbXsT9eVaUIBR8z9vtqH/E5lTcky+Qid9pai6zT
SZvTfwv32Ob0exgS+4ltn563YPngyVthU9RoH5ljXk1KP3/mORhyp2cXblP2Tqn9
rc7bhdwk2O27iAnMO5bL3jJwdcg+aq0b/k0tFCQh/dSbLChG4UtCmvhvl8NY/bkJ
ngwlteNwGoot14WJZpzbN3mW8uWYazPcCjc9Ou1mIjHXnGUi1yUXV4+mRtujbyGG
M2oXMOhsnKqjuBckGfpnPH1d3+7fLh6bvWKPQRXvMIcudK6ssq0M35w8eJ57Wpzi
5rjYau5JPMtd4i6mt2SKeOX22XHqzl2QTj1OaQ6CmJP54IaPhgHzL05Rqde8tK7o
HsbPZtvI07h1jN97uCajZOTC/k9aotFixWENHlc2VmrtSWYakZVZA3JqXXfLpo/q
IUacPMbLzVvf5eF2ZkHn04hWs6mP3rmVXuNBdcoLUVsl2MJQRE1pJUCIhVtF7uZy
qc5gmVqlwbZPIs1I8GSy2TRhU0Zxh1BuPSV8us8wmdJJtbgJPcFcrWSUZHL/tvy5
ANuKnuU4KBYS5S1B1lkJEfvrCBnts2KBq9D5ezXuJm2HQXNo3tJhk2adH3qEI5hk
j5IhqAhNAFvAf6ccKQdXTBv5gpQs5kAhG8/s1bkIgA7m9919xWzWZj+BJbPIW1ex
d+6iWbYAqDneV/07tLzwOpJCYSW5No+7TRf1TtFhJraMUTwdiQOTDUG0a1GxhK3w
sCughHT5aNGkfE/O0Gr/OgkdzFBbYfwDgkUuEJ1bqwHARXI9X2mvHNzJPo5fjHxl
E2RsIjRATrK04QKCE45PqSfazAQGkg/viXW+7GQPMTjGpjtoGjXZr1MRqhIKQhMf
JCb3egJhA2k/dmwryinqGFeGs7ZwScWKqGCUTWHOK5kJ3pWxKSRsTdgblODS7DdQ
HOGFW96VmHWlP7vHPnPBz+lJnrvccWv7L7jsaANlp8ugil95cr8jrAoFRY2SeCIk
KJ2efCkmDiIrPlpPJV3Zcjcpui4QVbRKZAuU1pNnKDjyQaKErTzCQTe62d5DrJC4
X/zpB0iA3WvBBZHSzx/ahPIVkRwlt54mlDLt3If+O6IhHd9eqWFFj8EQr7sUaxjn
Ep4Irh4XKd6W/nQmeSmZdUAstYXgy4S9Szw4UF58GojHArwCg8M+hLrCmlufWNdE
L7lpRz5671fFU+XJUP/CQ0+3Pd5Qdf8Xkik/7Xpqkgjo9qauOgoVoR0SBz0VFdn7
HIbi49//umkWIsPG1pzaUu3TVDRkmuxTXDYOhVzDsjm09cSpx8G/T/R5gD1V7FFG
3YLFTMTLm1a0eJ6NynH04tqBuqRhx8AfwsZm8VWg21E7oo2lZAUr60GLxuTuNLT6
yeiVYf+V3UEzJuFwi0GiFUIzT9qWvfThlrmD3x70lmsu3WYGZpP23wmLygP9skQW
lsxucfDEbzHvPJUUTzd9t/R/bOW3uWtcWDzcY6isBHZ3hhhJRIYd6zhAd1wqn+il
HmTnMemB79b+SIdaR8vGFQCKCOSvAHuRGuGbwQ4O/37dZ0uh4TxGL5KH96WfUhY9
cn7vYWZrFDQ65nWoovG4zDHDGCKBA0+8S5KXBUYFxjCYCngtu6hL3CMmlai7fEr3
fkcApjuy++yy+5AvPrTgMUvBS998aLZHjdPf/i5vpHC6AzgnoWxOfkgfeTBS1+vG
6IjNjodpSMbOPslYwoi2Lxr5xxs5y2C9CzXTEPkN9wUAOGUduCckWlXuUNZYpSR1
9oDYZUwbJW1TCw58BucSp8BjxCuPSNa2X/UR1xz6t5b4mfHBm8aWAUq+U2cyPbMI
ZSoA03kJNUx/2oTIKRyC4bdMrec5tZ+q0bG0GeZ597AD1+LV/9iKMuWY1Kjn4F4H
RECEgZ4Qwcenyp+v6lT2u/34KjKF5n89fA1JfQYCJOF7rQp4PROYDNgfa3HWiM4l
+6CjhK4I/fjPnBlVqFy8oQurOE6ypTaH7gl/OlLQv3CyMh+HJHEya+OIMJD6YJao
4HouKgKwqy0SNxknlNUycEUB78u7VZ1kI1iJEmasCKMox1XJHAEWb+IVSrvy1UbX
VvXftRTfJc6M0cH3sCdR4WhJI41FJnMTCy3F5cXchHyXKXPgo1Em0Pj2eRPz6YEb
e1pYkagUg7X/iuxzKhnWEV5CENDZ9H4fGDE304KHUqTTbIn0oVvXPfEAKpLeViAv
N75QKuzJ2x4kgi7XHnCTBVu3Th7+VaDtZ+q2LpvoUoeru0y3eO4dwpXmsPXmrsQS
Iv0nmOc2rt32TUSPT4fyzNlr1KtYQMWFjOPeya9qnTjlmueuRe81inmklh2DBF65
RgZ21dwOykyMosfhUZWT8NovGi4NN40satrkvh/L0PA98lHB8PTW5hisfaByMwFK
YWd+d61M44W+aSXmCqw+LjEv7ve+yx2oTpKQ6HZzRp7wA8Mg/vPBDRSOWEf/qL58
kIga3a/rUDBOTCLSA49GGPom63ZG1PTwco71CrUiL/FydAdhz5INHpu3YoJ8zM/h
4CZ+E7z60D1r4WKa5u00ZvjOxcHhkboQaEGI8djzwf2A6lTgZrJDIvkuZrsQUB41
qIJZXepfIVDH/uNmuEIoVDAUSywgHQqlvJ7qNVinC0mEDR26j4cbK8ddVuNC9keq
U5LhI0BiKjKraf4t84SpYYVzfxlMhxMhjE1B8dTWp1OWRXyLbT/tDZftRG7SDtk0
E7Ay1erCbznqzCGDYB47Kupo+woJjpMY1yQjO/pHk2sM9Bm9+6igaoXdo20QII+n
1HzBHkh2LwUhO0otz4uyzgDrbVUyj+oPL+DM9W0SW3oY2tFPm3KaUoOujZo70+m4
tpZtMQyhbhUdgK+8AAkZtASL++5ecjB949yAkxfHSi0mFe0MRHpTm6fFU6lxH2yh
aOGglLAEJsN8kmVwqJRwhy7GOQ108X26WO3ghITRJ1NhlDl6XErX3z5pG3QWAPg9
gAcQ4O7MIq3Vo3KD4fb5GGUA6dVF+nX7k3dvzouWkoFGuCdhmm9lMYdTwYKGomeZ
Q0AXchvYHXd60HDHz1eT4uEQDCHqx8mCXDNjMhT4ePudy4npax7Z5GilyMHrOYnt
cora27SR8P3cArJrOMc7rmG4zluFJpfTH4gycX5ZvfMcPFOvDJ62Olto6vfcllnc
HkOzA/NSzgeCHfZNp/KlG6Qs7hqyXnuKjejELz/li0NncXGpmtIo1IwJdEMCYe80
1lq01J28F6IUDksjAzq/Jk24TM5QQlDDXluedvVS8V5qMeukbNfsQS4OTpKgtjQs
mqWWtRHnawDl2j1dqLOcA3BsnTBewRYqvKmxxmpOFS3WbIyTRFBN3u80EFne2B8p
bfcIa5h2yXZ9i6Hw1O7eJ5zsYfj14YzjgllunDl4NOq4evCuNsfa08WKxAvolzCI
8HDC5GbUgr46F8l+GT2hKGXOeNQ0EYhZ0yE0SKYPsMMJA2CCjcKhzo3lptEcdGJH
xJhaLMME/mjUjh7IaDIYHrdkalB1TNUOdYsBqX7zgyBeUeYYLNhBYQmtObsCSFT1
p7NpmV0V+t1z/C7Oi8yQbu91egQm9On/hPPGPPEG+ZprCwnMQN4QwuOV3Y0xcSoT
mZFkJ2yhXeUok86SGhdx5zDRvlBv0suj/bOpdFY2TqoYwdE3ZIDY1r5Ndo+l6Bfs
+yaKKxpLuhF38on7//O0uYPzd658jjqAwovMow7Xcvpy7ONVyAkR9mMruTuJdomT
CU8CLUFCNxQsqmVEBuzlRdiO5mPMzFRz3hixq8KkBV8TlY0xUAPwR1AAlkuWXExu
g9CWNv5G/dtBYKkwxZVHZPdAOS5HRO5DMde91uwfmNOjqLInAoVmJ8ecvNu+LxJq
FiKbdTSynMsCCqgDIvl+44t7S7xMHLhTzfXJ1vacu9JcanWUx8NLdZLgt2IBL2WN
QuWOJXv61x0Ql20r8Q0ixzVKZYKpbOEVOyAIZ+3nvpNUdgSdrtm9LgcUAptAIuGX
xWWIbvNsr9OKvvHgpyFAdrhKzZ5NK0jiOYAKOCPEOKFBfIx6Vmo383piXNgOfODi
vN1yFXQGHBP5m7vhXHskWMKUwamdfH8iVHccudC1cAGW7CwzLeeHwOJv3LD+aNMy
Z036CBB8w3DvkwSNHUNSt0VvzZMJ8/06oQ/GXZ5tUyNWoZ7SrM9TNiFH0ztM9jBx
s0H1Tk9LHmv8bOxe9JoXTxqVpRHgOwkQeoy7uPRkApBpFxIh1NIBiSMB1ue42vm7
YkYhdGJk13id6XlkzT8QaD1vIr4tjUiMaHLi+80Gs4yq8sLqqPb0kIuvQMDyZpjh
ADmlLNBgti9nBl+ztoFQpLFwVOoo8Fti7aOou9q1Ldd90L5e26eCbr3FL7cbXEzO
cczzCH6Z/q8mOOP8MLlENwKVZMxNJVH2fxt3IqLfvXIBnmYexornowEIY1Cp69IU
t/iry/uv0Ut8njBzsM6T1XE0ivXRFONBSoCBaKck40YgVySYvu1N+DDIvjQH9qWK
TlsG0OfHc/BXci81t+N2xyk4GdtBquIAhpx1DkTHVRESp2hIhE3jKw+YSNlSXD++
kX40yXPj9q6T2kAf9/zXENE982E0tdlesrzGqwJpZZvZjviMd4VBeii7sVnjUTCM
C1cQxS6Sqgw0CwlT0v/uLz8HkSVsd5w3fnrFPy08zYDSs7XpbmbmRjaLnD+SnOB6
S5u+iTRoc3VtBVmJHa0NeNDWVr9qZru8ijrt7QKY7ruoWG9G6I1qTlKSprCvP1ki
fwkAiUKRTv2zXUV6qIpqd5XbkHg3wqcZFy3jLk/aE9XgH/NIASMF6EDg8S58WKBB
HhvZBYHZccI/DvpwP5X7F0hUDev1fv8gE6uECnVLJZXxNs8l9+l1WW9H704kkiOn
UDHgOKi20DpRs96Q9mG4lfzuVnofjbPbEEOzuJ6JiYtTnzMVwn75nAt0CbH4AIEX
sq35VB0BNi4AHGhqcHTGwhGV+JDPF4EAVwwJJNQVW1v0Bg2c4mtebycOmEaHIxxP
OTUcuirNlAXEXsUFX0AecCkxlbRB7Rx4qpEAfIwQxXKFK89XG1qtoy2SLvBpJ8WF
QiBIxgfF7j5qTL9bZSPLsRaIHLxlhovG/0e4VU7WrIjNmQ9hJ194HoiXxUp+c6te
6r96+CuX/JFKy66eEUoIULTG3Q/j+3cIDSgNDDtI6Ilm5WQ5zyrdLlt9QD4ni+5b
TNfoaUaPJNyATnLviaDFcQ8IEe9sQpk32mE+3A2fHdXWFvL9/mrArMBbsTkO28IZ
HezaWygQSqSdmN5D7e2Lt8G3rvrED66TzEXMzYTQal9rbx7jT1g6P2QuNT5W6EQ0
QhIkPr1HKy6Boyrb+b/JMaj1HVoS4HhAL6QJUOP7ZbIGiJemzBYdQ6cIFEKqfTH0
oIl1Vicm0W6xPKfIu/ZSxFiYnhsc/dMHELV3tajSMBd5/3L147NbryUPdt04kVMb
3JXeO26cmJm5WQ2TSkqB/PZcUUigtrmw2mZAulwRgjWP1Pz/coUHLfysWbXTkz+8
amnGrJTYXckD+0/C6JQqcUiO027TAFLpYelsJWL1miws7sMLHmV7fvKH7LpKPLeO
Ks3W8E4/u5pTSxpC2//Ptbi8evXTelQkZ3PneukMl1DblzTN7RLgNcZaO2rsTXdS
sCKD6F4q9ca129s0tU+OjjFuCxqBCKd02L9IyGJNbvrW672ZQ5BWb0SkZ3VyWTHM
uAtd1Gn1QDM7sIvdso3OfnTN/1V1Qq4PhVV+JvNRAFOscxpormn3kb+l6wDzXtNS
4fMsclu3FC1z4iGwkNbXqnxsuGgH/iAk1jMLhho5Z2Q0Huw9dJbyAOV58YzFPvge
5xEMNxYIU1+YQTAslGfpUb2C8GsTpISOQkZKeUoiL/k+/SgOiB/0jvI6hWNT0hOM
E22PXwVGhZF5swi7LZgzIs+0WHn/twz3izVn50STJY5CASHe8jU+I6Xygic/iMQm
8uYpws+/gbdYXxHWas9pDrNBpkE9vjBa19qj9Se6nQ3P4lNgjJrEd1NkyTNL9e3+
QpZM7nZBbAQ0qtGq+DM6Rj1Bu8abPsCZQaU/FjX1tQQR5a9gC+FbabahLe2+eJFB
9wL0nqtng+eWvgIvkmMzPwA3qG3n9oSlQQQkDgpTHDd5XtgzYdEX3Irwo/t2fQLB
V7Z0iPZpUm41BSZ8zb2b7HTyHvhr4xevS77CfNCyyTbmM5fAJuEiKq1rUpMCn4JZ
4iDc85T6SIIRivkXKVhUiSvp9NU9RAW2X+xMzcwcS9zKPggskL/SMtd96vFT4n6P
uk7A3uW9t6Zj4+x09zivCevDQuBPTOdPiBWaq0CyPpK7ZznvUgrM4ItNXKYSkRvX
sRdSYSflOMRjc+0aEnvKJVTiizaWvTG7SVcOudZcb4kw+Y6s94FcdBDR3YiDHjWL
pkE5MoKRpMoeKyfML70KAQsQK9Py0FGj3ypZFwsVStCGUjux+8j5yHLartf+BEC2
ITWSK5Q7wQcXVXxdWu26cV1n2sIsRwo9EllzzfdavzG7LMK7lHSghzSINLFzh59D
7N6xOqjiMT/SMGXU5k8x0tNDc2j7FCDeoIuM/Vt50crVyOBFAB2vXZtVtPoTKmpI
iXZhlLbMWKKme4AoN0dBQB9QQXE0korQj3RCQ2iHtH5sKY/OWF82XCMa0+r+H9GQ
8s3Z7wIVP55E1uf2MR9jfle3UfmgJdAH3Z2zwffRcfeTp6r/Rj8x+nfeHWs5m4Ou
DA4GT4pyayfVSQqKxyBKhfQlzOtwjj1qYBk9MbU4ieO+7AMNEKprZM9p1pPfEsq4
x52FdCSjfnkI7E2rcIxDJzon0Nhv3HBrJn/nxVL4HtZu7l38cGBP6+aj7gKSEmzf
s59caXFsr0NUjHrzhesJYYQ8PIsIH2h83uZnPYthAL6pdwTUnxrgeoTIGnaJ3gI9
xjPngC0F4NVKSc+8k3XrUDKJ1BpNg/XYdCC9FgPAFXgTOgdMJDbO79sbmovYqfve
es7N1tBSWhbAYXxEQY25pviRJJBq4nc8FGSAvfn3Z8ONuZRACb6BMgxXB+cj9I8b
ocWVjACM3527sJSh6cw9GwH94lnVTXLMLNiCbi+pWN05Tc91FBiqT5AYWBaPI4cM
Om7dROScuchYRydFfxp6huZd5HufUy5I23ilE8lyQFd33F5uPOQKbpn4p4+imzlN
62XZIBjVwJFWbM7M1HMC6NUQq10ngGyDhx/PN7OgaWZ8j5sAgj8CxDtDWuywob32
PADQm20rc7UtjIdeNd+EaGQzE3jtmDOk6ovFzyMB4LW4nt3WLIiBiFAyNekP7hXZ
qp4FVbg8GiVLwVk/P9CXMVbOKO1HX89UaGfG0+fubzmDtLsTtbZlN1nFyFfx9F/K
FujiZAj/0RA94f7kvhlVINXR1UEw10JBKZEq0z8qxFWBl7EV3AkivsqPFeNWdetB
L9lPtE/NYSqiNTxxbe9ZNMIp+Z9i2pelQaJ2RURndf40DOx6L5G4eYUpzL0CSSbu
DlQKvaRImucctVeuk3vDoSfdJIfIWd4NQRx4SYr9vVCcXKPBn9gQZFYv58+vFCEl
f7QAYdQc1eTP3A05JxF9yguGxeZr9Ad3yfLQt+qsJBrx9+WQ4rTOZ3hq1GnL7rfm
EiWiwiFAeR7XtdnEibN+BtfEhJfzgC/28OVEvw7pXEEc4ycOXw+sJZHz/RVRk70k
9upS0NUi8qPuTelu3Ru7hJ/lxB+yCDxtNt1UdpEtIi+s7vj51k04knu/EzM67wMg
ZSCGlGXTsJUZakGl1QPmp5t23mFBUt989XuOD8/CBLXBtxEF02G0whZHVOCwlv34
utfZbGel7pS32xsD9AoIJfIdoaPnklDPY1OdPchKGpcopcjz5CSQzTkD/BGMaV0+
TQcDztCQkxDFKGpfj1eoQ2mgerHEzusZ2nH/hsYybVbQZlZQX31UavrjTseD5nGD
kABPa8CcwiWte4Lu+dSSNrpA7xNPbeESmRuqeqAQy/n/pzFgUDTc+gdt/Mgnlfhk
3zgzcM56MPH1I2tMEmtJeCzmrgYn0EHwMS0hy4tNktWoaHodvU2JwcZM0PIGjJNQ
RVFo36OlQ2ynnsAnaeiRIfmN4e2jGcrCl0q2I9RxqG23wFGWCK9xqOPDg3uDXVVK
oW2hO60Nj7ZTgEQ+sIe06KISXZn+0n1xEDgeQb1opPY45ngDfuKfKeOx1CBDkgdM
8aUPGWazr8D4b5dn6Qh0FWEP30UXnLl3X8gCKx8dvRMcSVQBLxcZCeazMmNTVUnS
/JrGoM6/WxeQkRPI5q8rAs38Lqw2oU3rWmBqUPdMFqiNI6gxY1eETAL8ATIapnzC
hpVCnFrW2VxuiG7T2dsSIyjWvR1urISjqJTXUDHWsXByahC73R1qnUFp4Wyfubi+
8lqAc9KuLjFXK9WLM4TEKWt+Zg4vlRcO6cOQFBqiA6euKaxqEhp7Y/y9aSzMZkuz
b2pzveryC1YhETAcxmJXjLldfaCVaCtanCqiWZg1ZuyzqugybdRHY6Equa8mWf1g
HYYNdv081DhAhOTOhZpVxHhZHxPZT/a8oXq4kCdY5ALO595t27m6AbECuCX2w8QW
8yX9weKAx9KgCdtGgwnUCsfD0sHTNklw/vesd0sox4D3GF6qVz7McLbBzWRP2Tk7
+G812i1w4PQetv1g+uFkq33G+VYKjq0amg10Yujn+exHtDZwRsGa/5udRitxmInd
zY7pKtFM8qdwjm8U3+/4RMN1rbrXBbJa5fBxH46Kvmf5HfpgrSRVlamsncoY39fc
/9PQqm6C3TgKV2wUrwiKCwpm2w/E5Z732OzfN2rcOQcrx7NO4cpehQC3eVFuLcY7
ey/WOE4N3LYpYsTS8+Glv6EKComnugL+CEQ+kXrZzLNOUakvXEguRRqQtAFNFFja
7ab61HRmEymYuww8zi4wn83QkLP2fvzbGvVbrpo727+4YXcAWL1DUidsFEqjxG0a
bP/MESwX8lPwG4F7fjQHqxQssxqvoDPP8ZJlPrFX79Rb9Lu5fPnSG+w6q8w14cBc
GP5Ww7Czh1zDHHtcG1Rf1MgAkFrW7WK2Iu+VeStERsEDYf50mzkJd6SM49o/mnv0
Uaaxk1uehgkNe1mCgATuk9xF8OLeCeUln+miAb7doJULxgqXh+kwIoqcxhxfw1Mt
J63A5f61nFyVakuIzP1r6bUuVbpBTOmnqRLgOSfjJKqBwg9nogJdF1cSnlZ12+2b
5SjnK0EeNR5jJ99SCGCsjyJwUoE+0VdoIzDLftJhtMW8fjptxDyxTKfcxaF4LLuZ
RKrXZmqFx2Dw0KYt+leGZwtxWDm8ToEUiYB9cKQgNRhHu0WA7T1K0RlXhelsu5mQ
Vf9Ns1wR3qkThP4LBfQHRI++Hy8OGGcvGMKCwSuWIY8NLwKOr/7rfiJhOnQ0xSWM
4dNlTCCoKSyytujx4UdmVS3bUv62XAAP4FDwwXf5tFlrbCCa9Z9Gg8YCWIbQWiHk
im5bNCXTlZnJfZHSNGZXPO2tegzwVuO55/kj+HTLeAvcGH3v5zsCdmGF9x2RTRG9
pkHZNgjVi0/8H4d0yGGm8l9mPWrUHXDA1DNrKvqLgVaw9bmxM7SrRNcoylxqmgZF
+kz+eTFZRjO+Aj3fGzHp5XR5kpQvXpbmW82qSim6EaOQjjBZCdg3NahL2ovrflu5
aK30O/XvLMIN8YnguXPsnJy3DgfjS2OvYqOm38V3G/VJHiYWEDR/N0mmIXmtlQDO
NItc/weFkxrbsfns4dDhbMG2qYiXbcFDlTj/bBlnJx226MvzPBwA2g+SAiDngv8d
o8hiXyrAqNXIOyctw3hwqoYUwarBdOxIsdcR6MD8ZG5wz5ySAZujOgsSdoDxNW4e
znBg09pAOxD90kSlC38mx9E3c7+fqjwJzD4OvvLZObEvQUpGH6+ts6VpVVwq0CW0
IpEg5GflIUoW94BjHFz/Hs1ovzlDVroE6r1HjejTmczyxP+RfGDgJy38eM1jkd98
ONc4Yo6sicLmIUz4HvM2kb1B0nEACB36a2cL91GSJtmcJ+NIWxxMmHoducvcCd13
Tn3Pd7uQLR56W9ewXhQ3Rfi+zEXKoZkMxwp9GuhQSubMYYykmHSBthgUHteDhbAD
1vKTABwA9+ccrr7RquP/1UZf1FvUHdwIES6OnJBsxzmIyU8LmgVdTz5KsfxlSvjy
iEBoAp3V+i36XLSjKxUml4OHpnJ/eSkV3HEKn6QjwUHWYI/Hn0/UxhKUTmWzogRc
OLTiSD4eG9ifLplioJlG5IIRy7rTz7x2SlvPGMemLmy/zBlkDyP4ES6jIc1Uq+q4
akmryAbPSoNpCoJCz6VL2xZ8x/Rg6zP724QpDuB9ASrcZc0oc269k93EwHlIAu7L
n8bmwpqncHh0tPviUk9AWA0VExqxSg/N59U0/IL/kW4rHvRxnxuAB9PJeb1uFw0v
rl7a9ocdQNGf6oASkhaydCOfXtMhDSRwlDSxM5wLJuBDfkkrgGalKyCdI7baMpN0
fHWOYyuoWANDM7+RB73F+YCT7BvvAY508nhflHxk9SEpRLPDnsVsCv2OfpW3aysz
XSWV16ZX7fct38/WAN+JGYk0hg3VQedmNjt6ka4aA1q/2LVLg2zCEBTXg2Lod9Kv
41ITSxJxxJxTT8ctCWohkydMYJGaXNXdrw1tInBeTHn/NL2LBOF213PC9gnJkNbC
6nWXSZu83+wXcMjoeE2sQ/mwwwctHEogJQLfS8sqVmAKTE5LZD4nYDAiqGNcpGRC
dzsET2dxRKL+zFja1Q8Q5AXjIcwTPL7A1Gv66ABngTDBsrQqQFrMM8gvrTDRAZWb
Lokw4arfubRWDLhwwTyBxFUtXdd6SlY4G2Gy4Luhrmi85rDwAaT7OfisAyIpoHen
39Oxn8pbn7/CfOzhrwd5GSogxvMYF5jSPWZMcl/rh2pBbpMOmI0fccSWGk6T6L17
HMuET8pDw5d+l+9i8nlNm7abVuFlxvMlcd7crqPsqwOLh0qiOHuQowhAIq0uZsQ7
6DDnBydJG7MlzwknbV2eznzdDgvl9Gd7qal5f0BuJFg8ULWDLh0McRWejoRiVHIW
O+mncmiAQjlm5sU+t6YBYSjb4O9J8yUi51g2voS5xCFbVQ1P2qEOceb2Dd1eR1SL
nJT5xfXaeab9cQVdpX6YVz+ytyTCll8yqHGSC10CmUavlXVXBMmPbJ7nxyqOyT0i
wBnkDCg4NLRZzNbhHLtfopuISL9/TKMDdo8kXc0fVn/Dl5gkvHeoogN86RQ8tO5/
u/8zB94ArM6FGyuaNyziQsWAraKVZDHzkbSgM54XCkOCtsU0Ph5nIohWSNOfezOk
fTiT+rrwq22KPp/9QL77btDPF22EXDHLJk9c+VjkLpuP4lyi2KsMo1X2M1V9f6iZ
AN6VvUVWSvlnOlGLbYVJf71eNwM8TyFuNVTbPjZeueaCMag3aRU/Q9TL06M6Dc/Z
U1RLr97tWboK0KiXzvD2FfAOoAkJU/J+8O0aL5nTk5DyJPVfgzzEyKZmPhvJhEYD
nnCnp8og7hEelGb+oEGpXz+1PiBynIvVXOzakyYkhCtpR5pojReAo6Mfk9FXCfuw
0Q2lUssIre3JpZRW4Ya/zjpFIcbHjZk45Q+65DjqHoXXDAgYc5VpYTvGgAiP8o/g
KDQUS4uXpro1ePMk5NzM8xY/S3IjiMuuribEFTr6XMi4Kz0ai5aR4DwiXUZiCoN4
eBB6L4bGhGOK7vNkg4OQI8JA9CCo0viBcMj+vCPY6jGYhNgQIHwXFJpjJiaUQ71O
Hcbbq0DeXyIc1uhuCVd1Q6Bw+d8t3Lj8A6vIwM5KeMy3aCneajws0WZtxQvQOKWx
trhokQRvxGBFWAbO47vn+RWnMCuEMdPe1DY+KoPflRQvGGKbi5JTSrmkzA/9/yW8
RRs2HkK+npwja3k4Y14f2D3QzZ/jxWfmmwcLcsvAUoQZWr6ky1UziTeuuqCrerDu
Vgc9bmD9txjoNa5W4LOd4BANXJX4lS4mpgRohIxtQI0ZKkCHPFGQCMocb4H9hUgc
1PgtE+R92b1d/qTqFvORYXLP4A7ofwG/RQvmoNbgrwcBipSMRSUr83Xb2Te32lfa
xlpLWrzEGUgVQEqF+eOvxjdyb/I+6PG2L/k3LalRK5b21LYmQzbFPBNFWGqjA/Zb
HoLUCHU3ICblt8z343SWKOQYy+lhSP2QYNttA42xd0RmeRCdvsZuzP2wXvYjS7n+
iPtdid/Pqsv+KU4ANd7XTyTNQhHPv3hu6GuChZUoQbN1gvBpcmhotPen/CC37sPe
F/CdGNKO+JFEpJ4QEXCCpADL9ExMCySoCZ/oLvzKnz25vZzyNJ9nJKOA6cN5i/fX
lROu76xbKp+WyeUQ3YdWPvwPSz9olnfl5/vx8Apu3agNCOLKywkRBu3El4LbHWCW
Tgi3PWYWUL3uEiVFYzvEM60oYMQ/aogOn+7p3oF/LwhrEg36oPfYwPnLazKGE8rL
Q2vvLb+1eu+UF++Ar8DwVIYBv/qBSuxIT3dwEVKNBUjYSra5gS+7OVXUTRRIYWh2
Mkwc540gGDQYH2wEb+pP6FCCG/aExUw7spC9wanSTuVbvaXe1PXgwVWMQ86et2ge
yAICAn5yuX2/K4y3SlGfSjT5FlHsOPHhalfHFAPZ/3nE6q88uyH3/6y9i7222a7/
elSiFYmg5RpdO9nRTusMTobWoKQDZTLZ7r1BfljPKUvs925+r6k99+CzdGUfTsNC
fVqihK2QiF7rb0YZ00k5l2kFon+ROq47zIynN9vQ8kt86ETHVB5RlwGE6+Dm5n2t
CnCEONmMb+djJ4Gy2kcTogyFk22xMOWBZs5sy6e1bsauC5hpBU9wXL8f+1yMMFMZ
TAhFQSbW4xA8T0lyecAdknBM76R2TAw/+KCTWNE2CKtm4V4yaLsPePt6dStoSGDr
5EvH/tmU2Onp2J0D3rbloeM5iSMwt4z5fiUoEynLaAEbq5IRhaMY8/lhxj0Z4T93
WjeTvfwD+IVfEuyXRYRtRvU7UFsR/QEO0cLmSDdO/8ylpTgThgEJYAbkr+yrHU1o
RdO5rqechzdmD3cQrE3hIbDLJOHL6dKJAnKwKiLyv2LktKVpZTuEVu3H9oZSJLmu
d5dEa2eioTSVh2omHZdrZr8LJ73tyWpO8Ccq1597i+DUr370vaeTWSX6T8zxbd3u
0dzd5skCJzF25e38MnyTZeCv9+akcMEjqH+XRWMsdKZ2sFmQFDBL8lLW5g5vebkD
+Xpdv0LtyW/l5T4HzLMMqT/qOGVDTi6aaid2mZ4k1GLGalrnBtnwP1M8A9AUnm4N
ytAlg33KdDoY1YLt4UT83OZ8zSzutWKE7j/L4xcK/0BLvcHww9FlZQaWr+2g5bNU
Nyxi/X3UwmRxFoF0QKzUhEydnmo+CFhGaykz241CCLAAeKPdQw9+hZfmXVZkg4g2
FRfFsd8PjXGSHYugwhuYHplFoxjOyJozjJrdRlRBoIgpluv5dLSTAyLvMszNnyZ+
KhdrHmoTWziIL/F7TctRCNYDD6abJdCDhE3dYdnNEym2FTdEodGHpOPP+UBS2Trw
TJkxdeMv/ojWsHOSOXa5Lep4mLa9T7qGN+VtW26xylcopkUeHTlo/wh8vdMN0gxX
hzAXpHQpDABEPbKsJxFYmuHjCNubs421XgKWA/YLM1vliFv+mOorvbuw9tFYhxPB
NpQ+u1gxiw/dYsO+U6m4rt3G1g4JcJl50ZmMes6QEBS4EQeKvRDZiKiqSFyoMupB
1mxQVcLDxoGDiW86le0yEJygvivNgZhELYe25lQm7q6zrFEf4hzSuYiXsWeZAZP+
T5WTTsnHznt8McUcf6FLXk38doUWacoFdMKwFf1zVyrmDxNRKbUkFISW3ZodekUf
4Vb7kWgGDNaDiraBYMirjN8wMzFpvzON+h/HrWGuV9+FHCEk8Y9pIbBzP1EnexMB
0cCwMYyCn2s8a8yyUHGOVJkvLRQHOlAlPnxtSzd6NG/uvtTqJhlrKqo4M+4lJKBT
LXdFBFxKfw3853FJQNJGF8KHCQzSp5sX4ClphiWGGAq650bn2i6UPqoQiIA8ynD2
qYmd1Fbpp9Y+EVI2uDK4p/y+CwC61cTcchHnjuwgvNAO9lRH/rw9BBw8XoJNs01r
jBAvhiCx5P0BVBS4kXDyJIMoclZoiPG74/voE3msTsJaSDf88O0HbsRkX0cvUotL
4C6SrGsicbRcf1G0HBpP6J9owUuqxl+RE16+8JgaghhEO2ETowgp1A2pzb+c2UdK
waRgJngJpi7htnzrpc8Oa/uJmADbSw+0dYuUeNCGCL+tBjW4qW6/cArD3a0VZQ/E
Xd9+FjEOx8i0cDyuWZqeGYzOaouyBOZ6tJQLjiJ3K9Y9nEEQvibiSPiIlbQTt8E6
lljKDExwR40S+EzsfXULdbMk4mfbWwYizbLQmv+8jZvLA4qkBhiac+lAVJECNZ7N
gnBmEQ6RR2vQx053jkxm/BpOUjn47vka/wxCLcl01Yc0Zgu4q6aesagJmNsYKvog
/k4DO9ff03mjLTtRsPebdZ7Y1RUHQnBTJNhvaZo11YAT69aheWyfHHaMbCYt5S8h
hO1oMyV9JMDPFa9B1YoXI4bmlIGjAdiUaXbzX4QhNDHcG3e9Km0hfeM3ZV84PBzm
Gl7WM8Z0AMNhTOh1tc6VOQNcMmVga9O3VNP3K/fm8MDry79RKiKFT7JExxCklO7B
qbVC5P48YDAbl9PBA3moaetwwaJLRk+WNu+DE5kxsPxL8oxKCsCf3XPuE+lBXaH7
HpkC1KmI73KTyMZ1AxKVvrAwdzGx5yGjh63hK09lgcSJLQh8xxBY1mFkN50xgCSA
vpNmPUgRuEbQOfBWDeFDx18k2VIDqgDcbH4B76puAJU6hv55j2U7cOmTswZ2Ez8t
MKoC1a5oVgkEiKy33gzQhGQTsfS2ptiARPhpr5Zea5dT8BOJ299f9JN4aJNiW1v+
QeS6emryU8/br3Ae86i3x4TLR66JWxFBTQun5XSON9DzoKLaBBcA8bZk8pSO0A8Y
sIk55CTAkVndXskm2VxukKDOzn4rCJRFLYY/ESTCdhWQhLNhpMY+gNF2QAVlyJ7H
Q9M7PyN2DUBEPOGI5u39NpJdJj20izSRokJtkrjYZcPs+Rxg9ejaPKa+p9PCTJ8R
mja6aDUtwMvunnTiOBAp2hjDAQzrkuuGtDnuAtNcCHJv4qMpsZ/n0CMjr+XLoK4q
Dw1trTmDfmPtNA1Va+3vryLP/lrfnbFxyJv4ZuYvKZOgpBs2X7S8K/udHlaplrGh
3dNhkK7yeTb5aK6zjAB/N9SmrEnMuFeUce7/sOsDAP1HNhXMSiWLTW3BfcHNo14G
u2K7tyZRK+7vhM5s8g2v6yDDjtPvC+4jTsbS+SRaKpd8PoGHFYmgiKdBXAgnvKkO
X3TfGiDabtX/1G+eOlHO41/qEoVg0zf7LU+MmOM8UUcpSzwG/f5iP1AitqobU748
nE76mZlg/Otw8yq9p9Hm1qA/h44vHZnC8/XzJMYo9k4GvfeaI7ML9SrPP5r2GBi4
yh6odOYuu99bUjgsB8DHT5zUGDnTun2NLwC9tOEM0WWxhLl4IjCsHIvBr7BzWXB8
VklWrnPlDSC7hHbQaMGOHRsdZSR9f6PBCeSxHddtV1mmgf9tFuUSr2wBIUP/08YH
wX8Jru0DYC2fJvUNcp4rmezjGkfK99n/kD1o2KONPiSvALL9GAWWKhb4D8FMKPmI
MKtRrqUq0/WBn/pr9DFVt/hfpAVnXGqaD9Z7C4atbCaxbFe0rTbJoaZgOdhrBiQu
8sUzzMX+me5KrCd/7F+Or0YZD0QDT0YWW4O0lkVlgHPBQlS9KvWOhKDBr3mxswDi
79x2hvKdaNTU9q8CA42RAEmSHUmmlbdTn/wIWaU4QZonU7UYWAagbwaiL+KvCf6Q
Ig5grCLhiJEjhVbKx+N//yror6s7TBKwNDHI8Ey2Gl7Wejx6NAOsSZlAHlfBUAt2
0EzCBqM1JSNASkuTCE+6GlB50ZQIWHWXmtSrOwQ37a/KSriE7JX1m9AKg+ov6JZ1
fVa4k7k0ydKrcUmTe8RPBUvAvrpDfOCN0BjzJHCrr3e4g9LPFhw9ylozcRnh+6ye
5+IwsWRkOr8xAJly0R/XxIRvRoE7diaVkSkpFCYPQ7k00XFzu4DvadELfv/m5Y7l
dN3cOjmaDJQ3YHCIC+RNXLhhX+EYpuDUhVnMumT9NOWtVkn7Jic+0iCsAig74jtv
JwQyEyNRay7m6ILa0ulivGbGE1a+Zuz+jTD9Ea8rb3Fd9X/5P4iA2mObL+PkpQSZ
1OC0yP9A7rL+MAzNCzSQxhtlV0pfYcZ5d0fu5ExnTCoIN5dQFNb9VNlKqGk40lWW
RJa6YdvLbKb0NKlAgm/Ysl+FA8ohhL9aeRoBZKTLYoNbeGJRC4DEAkww+t7n9yaJ
rEAv1C+qcTAWHftRdJnxzCfEfpB7CLU3RF8qCK/DxAAoxs5M3i8ny+tr57rWVzmM
E2wowkx9PzkRIth8D9csHGnQuz/BnEtHtVE7rvW6BUZjNvGpbGmBQnxXPGlITrA5
XYbB3/khHyd3ppE+6TJvNOAQIoFLp31Lfvv/vvatpMd2L2CS2I6Ut4QJo7UZoT1S
PHU4IiinDXsiXAtbEhLuG7nH6t3Kk7rfKDQ8AOrcIF6XmXcPrdXPIyxAsi0LMgX5
UCP8GYWkNZEZBeX3t8TypF795sI/TwaeQzIe0o9TR2b9omhgb7BuMNV2fLceNVuZ
J4/gAlhvCgsNflkd+awgointGp5HGN4Cz150HA/+PQTk4Zm8PVptGaD8+uzBoKvA
eTG+xMMFH5wBQfT89m0I5HGRlzgRbuqduWYN4uXdmFpWUmNslid1XH6+GTnDOE6S
UmET4oI4RypPCDXZGJDem3gTTIw/nCLRHXfV8NxL0q69PsdmVzpZ8w3OgMSv7yQa
ar1WVrL+MRgD3RQvb2yRLJ94jzBjO2UxRwkzAJSmqjtIQTYGKuE1lLqM7wL+uOhH
bJaYsl9IvNl6aHz146JMa/Php3QflzAqol0wZ12G3aQURymDT/h/Nd27wNcAzofN
2BjEdzO0jybzlcocFvThLFXXMp83RaWExY+73sZNxAmXNvUyGnMXewML/MN6OXJj
fUmxsqv6DaisMnjXycmUcEsE19NzKdBZojHVM1skYZ6udO43zIGE8mI+F/WaYOu5
AspYBnOLv61YCgjNCAEaOJYlVE1QNGkBTQ9RSuUaIFbdqDzObfBuXmOcI/GzMYUg
X/plfuqFVHWjF7MPI5RMMsxmrw9LFEjM3vXyH9XTk9r2naMZBd4qgXHUTnxZ73cn
Ndq53BRukWbDCEORxwy9x2BSqOEiEqRZkZUU7ujgY6jMZOnFOx33cFqiH3Zfk5Ev
2V5k7ffxPY3hI2djaY5GfM1F5iAGQ5xVDx/enVyyOXMI5FhYlTJgBLBDSWeYSBDi
hdUAYAco0vN/8LN4tI0iM9PJt88OtsE2v+BPB4KoKkL4e3MHxL5NI30LBy9gb5AD
yiB4G0P7ET/TTOVFJIYQxnhd9pUDU4ukcHVAVunbMhUg1uRFDqGBR7HIA35CO56R
oj5vOrMRcrncnrVso8hDMRc2rVFJSLpQP8CtgVNvi9qzgZ0HDjXMjKi3rISppzts
2i1+42ZCsKTy0aLh0RMT/Wj77kDF0IzZ2dBHutF4f2VCacULdXyfKVuYf/3YmV8H
9FLdOACPkmMiEyGVjvOMSBjIFTWAYiAv3HI0+DMRYPJgocpzCRjAExcwaLf6smfM
7JtVT5ZAcndgtRXtRxunOJcN3G8jS+rWKvNMsL5180UHxuVygmTwCJyMFzAaMShX
8pFUki9IjtLE88xYmgHKToFWonLbUJO78Lwvgdp3vXRPT1tKpj6wbgrKjoJJez7V
7gaZ514uidgsn5SjdibEd9/lhyuabTQC5a0i09qfkNHrIKidFx8ztqSF8ftlxbvs
hEwPsWUsrfD3GTBc86ty2UbhBjL133pDI/EwlYv7OKGnkNmEWj8emAa8/8r3nFJq
EgSRntI0HFOGTllwk3hB7TEm0Fi7Ffa89DbLFQclDRYrSIBDVn8wwxsXhCmmvA5N
EHQIKKqcCDQitV693PQs4BrQaQtsW7a7K2OsZ0oUt9JnljYCuJKsX0Q4Fp40PcV8
80A/x5nJCqzxj2o7DYxUQYSIvLCj1ZnIPV+NVK9gMGyjRrAVpiO8n307KSWxKS41
6xRR4bS6lQvSuz+dGocIm0fzOHWLj5vWdYL/VlC/QMFhQ5edA1dLw3zk3xqP+Crc
5FF0wf4JD6MGovznb3XICwG77NyUQn4XC4AITd2xVkBBW2mN11u5XUHTWumSnp8z
OveXNMLR6kKkar4d4tciA0T9ExToDOq6KCIB4y8tsUf0FDvx0sR8l1tc31IiLxHK
9f+8fkdrEXcq/bzZzKCYKWBVxYVnCCb74iqMTgu2DA/yZcpdK/QEIokTT+aNHKLa
xOHiaCBUaIhvoFUH+CM8CV/j67XH0UEtOPkknuV/NOXUe44avwp1bByFXqqQyN4M
QUVVNi/K1NuvMRkzZLYONkoChzRRJReAvffm27xlUXbyVnOIxHd3eL+YnygahsnE
hpzBS4Fo1jbZY50mr1xhkr9EOjJs7P3YdI/dO1Z1q2Sl9eZp5FieowWp9U+VsY2i
yNn9EH+l7u+m086txL31eU25N6zGtru6IZ3efe1bPyUiUziMUPrXy0UB6oJwfUXm
Dl/ASq2WipgXMxDWEajd3ZM0hcKqc2wVcvU1OOlcdiYU3POg6cv2IfEFDj+L/Bip
8BBBB3h2YoH/2iPMI/x1W8386aKR+zzDiI6aLyltEX5vBnChZvGvnnikIBPyxkPl
6rnS+LKEZv/6OP7BN9pLYQhv0WxpuOhcZCaGojd3KpQD5OG9UsStwOKOLBW5ORKy
AeEa+c0xIbMrxWBjS8H9rKy7qZXMoYbLY4/Aft7St0VLYbcHT2XoEvkMd123AWt0
wtrPeGdTbHtlG9evpbb0hsvVWlyRfwP6bha74fq10NA7YaDHqdfSl+g6NBvHf22l
mpzlBMPGC7fzgnCJh8KoAs7YutNn0kAZ4bhx6G6qAd6fsy32fMtPxqFb3JA22Dzx
mzJwO557gR1q69/eZ2GKA9FLD6Z4KNtqugJDkXQVVdqTyVTn5ulh5o8aThECUzY0
wxBkMVTYCn8rj5kocBtutlFyT1lX2Kd2pQulsGETa7c57RAGwDcfcHRw1GkP+D3E
JK3RURDZchyCjv+oIoafK1MVNtweaJ0nzUpkaQF4AuxNsY6heXSqNCBWVmx55Muj
O0HLoDJQ4u8QwyPs4OQnhiPFpGveWFZ2UUemeaHrjJ77uIvgxsFHwTyptdWxbwCc
CaQlTDdvA2vlZToTTavBL32yEAQOqAR8JiTmUY+i7cnr39CS6ed6ImE+xzRVfAfi
ofS8ycWCm7X3R5nJMwLkuxHeKi47xZQ95kqyR8GvUSmRE3tlnVi2hk9oPkGBaYB3
BnWzScaIja3TmPbrCG+QlpK0Cv1/Mjq+u6cu6Ufj/dTRVGkA1Ib/VmDrLx3ZxRhG
xFkVcBX4SQ7nJ8Oq5CcN0a4f3BTlLPWUeTHyBdbhhqka+JdxMJy6uZQzp0APKCB8
RqyjgC87IT1hrGl0se4GRNo9hUSiezQcTbVAXL42AeW3Or5OJ5rzP3jzAEhRM4iz
Sbi+fDqnzm3IvF85LkOqND0e1Q2kUIMDrJNV6QzfM7raxOPTe6dqNNtUnclBkelK
HUAMxpe1kO5WjjuLNmamcDoouVLthML0mQe7xhVUXuKiaWxaRL0HqSbSolUiVygA
17SdkD7i+ZdAssIZeMfeKfRD2kapa1shXhc1hVeDnQGHlEuNhynaGno6I09rY4tq
9avGVD9fYZyOG5h9pgsp0V9Qc0rg29clda77gaO55cH36wZKGkE1OX7Zp+CMyVsL
ukSy2AyLtmwfEs99FxAlg3ZBFEmSMYMZpBSurd0EEZt2gxmjCmnnwF3xOQSxa/pp
vYO7Nnorj9sMEF+m9Q5LhRSfaIrwBBSGwEufgOUgmM2PtrFzfpT7pI/ZHIIZq6Uz
mcUPMGQY3uzq+F52Rj1SieLoj7XKINp3gUu/+pF51zq00SsdGblqkGFnMNBqCftm
4IbzduuQ8UdlEI1UxGGShTOvo1nVC0QSKyvW/+VrokGSROddj1U8vfuu9CBvWKmi
BiAUIRreiFr+lHFfcp+JHNS7G7Jrc6d6rO30SppgwVw+ctSOC+X7lA8o7Rjj0+8s
wiBmOTdyjP0i1qcvOeqYtPhrAZ1+eoaR6Oyakm8NK+2MWQGsvbAD6bIIsaLdMaTb
zLh+wE2/5Uyf6toD+YZp8HPDN78Hwj1y7hKbYyZPhy+zzumINZ/zCWLWLkn37oI3
kIvinv86CHht9EX7h7RuVAgGo8rN4fzGwpudpIw6XMetIeYNB5+9PZfnCBCLSH18
oOpMJanse19TbX7AC0qS/z6xjVJ5Ym+gZxYSfhgpSJI5DWHdZSz3S1z8sEc70asX
xh1PSKnv/HIrbBxCZm2KN5Q1CPhsnYsoBEi3FZJDTv+ij4+dGzFVmMBXEEh1ozhW
1VwNf9oZustibbIhJMYZE0PffwU3WtV1hSLIu+aH3DbJBJlg0vbPm+d2ri7DqM1n
r/bCnb9wMvJhR1qyXRp/aa+h8O+CwFE74FMzFK4EVMttyq2kSrxa8yhT7/FgnQSi
bvylnDXuylxVwcseXaWV8Q5X62KieKkX8biw79hnNwJZFCdW3DJB1y/UREaVdpH3
KfW0Ssp1P/MRCTTbjGDK7O2tcObf9EBw3r/GRIxxK2IPy9W71AcWY3Gogc3xGXAf
tHvZKudt0zyz9uboP3oYLbD1oxzWQCFBkJzlv0d6jZ99awxW06FaakTIvDOjWA+w
NixBPI3Efu3GTm2qM8ZkRXNd1jMKeViDGIEhtDnIUzL39ujF8xd5zpoqNwLhr8xs
Rkin76Hgj6yg1C2PDd+dC0t9mxZm4VpLjF/tl3lg5Lc4QokBDSUiwBRP1qLgJk1u
pfHye/x5PAXuxy/tsY6RDMQliLg8HrQOOfqdtiqOQBX1IOtR3AGNoK09RS6yKZxk
V5HIuhTHxYkKqSYBC8uflhBqDFhYz0Il+JhsQPX597BjDG4NVixBVbEH7byg28lq
myw7bBq4nTaqXIOBwsJMZUDqfiqDkeDvmbwEvXmHYw7sxJDyTZnFyXPKdZ0aUc0z
wyr+LvviDHfAI1nEyBifZuBaDHA5aiXP/AVxQ/OemM4dkTKpg/fl6NYHMF/HbHU7
+PowTBN/5v7uMsk2O0yMTcVK14R5TLtkWmVvJzMfuZQpruJiunkIMCfraWCN7uSG
0+3aNchVH+x4LtOTCKTAykay2kw3fpMINlHcBc0OlHwX4r8dc4nLSP9xBdG1Kiol
90f2FzJ2FzY2Ubs28fZrIyVbZPjWcwOP8gZz13Piotyg7Dr6zUefj6YR2OzJdQ9N
2nU8ELIS7EXcYD+coicRPgcnQkVGuzxETgbytnJSKtCfrjCxtIjaXWTzsWwGw7NO
3uwzNaRxMSSM2B0GCNgfRWwRQEqhz4QkCmZKpTbsGbOOGGUJXC49DNTqpQ6C+zBz
6hLY5Gm3dEHZ4UIwj9aA4Svc0Rmtv6y6BTKxxM2b3Dnt6pcVOhZlRkCP2y6xlcuR
lI8tt752BE3T5LMyWYoNzx/8pv2n6dPWgR80Lx9bfhvj0nidq+JC5n5LirGnsaWn
7TMUY/ovmfJqnEmqPNW6NJt00eHisrHmX0rre8/namEwOobvpHgLyRH7yLonUOaX
Ex1Egbi/yhpvA2u4b5bTVxdkoX3FeWFf6q9c15rMHF2m72ER/Z+ivxTRyBx7vCaC
ztR3mRt9opdIYqTcPjrq1EqoocfzDwgMQ+brCXAf22HgzfafP1zVy5hhWGyNs/sx
JsunD0s6trpaG5qPz5kp/Q7OvPwnYI8YI3TEGXn4h/hy9cUIIsdO5cSSdeXsbCsJ
orOlzY1z5BVmgjPJ349B0sIcYbT2VIbOAgK7i1kRaGmd7BiFUmv8PX+CON4MGgNf
BPhGHtCmvlLR+ph8fOzdUzfY1f0u3sOF/jgypOTtYSMGXGnzYFmA8HWQUMFHET8L
zDoQcOlbf63CfUqTMlLzhAT45PHkB6UdF/EzyBbLT1gBKuJP0FAb0dOu/e7mIHXd
2QFSW90k/G5G6y2OLVe4rAt69VVFz3eZN45JB5EhqPQi2VG83KzTXQbuKDXxEO3Y
Y7U99aya+ZufOKgyCX2ZJFkkLIfXxAxGoEjDB3sjvEPYWBi5nmacxPlNbQSBnxZ6
xZtPp7Uvxwfw3PKQQXMxmgfURGIiasaqkPQeQzzcb+k++fikB21THhOrmnlto+O9
Aggno+o/sqBH0O5VdqsZQg9Qi55piDbFANkvvIlJEMNDowbvtJ137yOn/hapEd3c
MlfkSdXXtsMYFxINSzCfq3CD8JEFE6AEGtoWeoOrD0IhFhyiuJnfA1EONmWVG1Nt
9v6UP14htx61Pbta+dApp7ioREnYH3SBMr8q2MHtNXOpb+PrVE47gXMbMwY5NeZ9
+0dC/qftTLQNUzqP53B7Nn0I2gDSRA0Ix3CIB0LpRQu68f2kaXoqxU33dSaR8YdO
Vs4z5XQMDWuGSyMnqzBwgzwSo6KJnbnBvXcPI+yt/XrtLi58KN426UaTBBxSUfwb
OErYbmC01d8gmPSQ//LNspgVM0Y/EmadJP6HA0pxf0Tv3+DVg/bYkhhDV6NgqDhe
PDz0dXA4SxUHxAkFnrjsGJyVkHjid+NsGqrwG+JBSIhljq1/k/OhLxieON8VySvg
28S29RoHO+GlbLoqPThzEqh24hTPGW7lmRspZJsyZOkR9NO2Rpyk628CbmUylJLY
1YqRSpiFDr2CKmqPwiMqkxg5Y0eqFbvc//qCzTx+L4xjz/NevSgDYeuJh5fyal5s
2AxbBgkp0Yy/MwpEuyYXksjKpG+j6K4qyQ7MFydRNEPvfPUHj7gwT0txhXcGzRbV
m6YSJCtu2WiEQOQcV+97tIYlKQ2tJ7OssjW7ZNOKVujT5XDXa+zG89C0c1QeJDKu
SKP5dfxROJ86u1QqEcZq8SvSErMHGlzPH+SRGL5R6I2SP9PxsZLKeqXqZrOBchMW
V002BwOfqF4/HsOplwWvxO3oWRjRmtF13d1SztdFIDlVJEzVdWU8TXudbYC+4uWm
Y9mMehrwAD6m/Kt5AZ5x4TK/+YqM8OVA45csozLlmJajHLF30CfX9DmqU2V7uPAl
hUEnk+IQq0+fwWAxI/YX7NAdKKm1clasbVShaeumRH8RQr14Sr4upvkUyh9UL/3l
b/tTcygBdHgUtrCUdDdgXuIc+hxrI4kTJ2TU2hyg+cEl7sOspoA91DVtMr2wIUNz
XpZu5Gs8gTWqkyUpHwTrmJQAYU4E11wSmwOefRzq6QDNp42l1W+N7PuyUZx7qy9N
vxx04R8bZcCfcYwy8A7NVzELeqvJ94sVmtFUheJYFyq2h1x2YK3j4dYz7ejk1bBZ
tNYDsswwD/IymXTP8vxxc1kDETNtehATnXCnLYjKuIHYPERtsCJjtKwOmk4BtnHR
bjeiD2/Xt+uQZggOpP03uaiBbWksLyMlPT7QOFGlUw8HuOlT2Gm2ZSWvISchLZvf
NyRh+bvAtbkpzbKvpVwKshE5agq55G17ER6mqdNYAgS65eDvyPVGJRr72TdAeq+s
AFiX0t8NWT3bRlayZ6UdZCbfTJc0LswGrhmOOAzrwJHiDfSO6eN/WNmuqcwNdniM
lM9XpZf8OEeyJGz5xLay5hAP+SUnSLbu5AdM1RIexpfvNxzeHq+l/y4jyxyZerSQ
2wQuCQ4bNZwLZgW90KoFnIpKlfTpAIgcFSjd0tp8e9yntBO5wXD3vvLeZDWgnmN/
X19YbrNxU1EeUVTaILHD+AFxvsxWze99Cv8C06fAM//0eznB0Cl8faJ2ETrQJ7jy
m5NpibrVCzfh84QaYzLfGH7xJerY8wi8ZcvPQesJ6c8l3xWGzJaShV19lIB1Y+5M
3AqhLP6yUpgki1v0vn0SQl2jw6f1II7gOZUykOFIx6GruDNOjmPaCSHVneZkF4xs
EaFiPcSIaIHa8FJJkMShZatHa9iuViHozc4eixvjC6EnDI4jpE/AxpG4+tXVlieu
wlDJYaf2n0KRXw6A+b8XeCOWYgKBhutNXZTV7RMhPtqt2279wD0Pra7MjToYJYLe
fEU/2CKCAmHaz2ds+drh2CrqF7kghdDroPQL5yxC8Ms6eeLJ7zH4H9BsRPWfOKtd
22Wy7+V7BykrgUrQZSI8aQZ/JGy21Y856XUcz0Nzv/eY5mkBOILF4ftbQFtQTjvK
6p/U/9Zyqt+WBZLwDA7dpiTmfUM6O3NKkt0acv+EhyOlpCxRbBKuwAHXU9X7Mv/4
SMzvjxXEL+R7ooZ0hHNzkc3iiMjd54OKD2OqnTkY7Nfwh1+eFreD4t0w32EmDSCq
wx82qimftSMl5ZqxG855J9QMplBHQH8+DnAesgH8XerFaABUgTF8UvRfWP876Cgv
iYlTvn9bsNET9tNQS4c7xHYeKkBrTYYOv0k53Y+CVBpXD67LoTDowa1dk/9/cIn9
Y7Bxc3B3ybw4OINV2ph3woq7A900EygZcr1JiIM+F8zQMXiS1HFMT3oQHFyLX5vT
JdQF37MCvpN+jMoK1eQCbDH5kvw1/HT0RE1cB0w6bKfrYrv5mUSBbeHhwLLJw6IT
TLbOCSu8Ta6SY6dsZvehaFhgMA23FXqvgpSb/iSo7yoUVV2OCCKLh1jI2cPm4ZBA
x3d1cKqSiwILNZUDS3UtnCgh51P3kLi2qVSnDxeWbk8SyCXxaq+tGFJGQl0Y6tUj
axeisZeHUTglJh2HbLr6dTnENERI4mLtNIa86MEBMWTPcUAdjbS7bWtQnqaAGu/W
yFI4mZ8wJTmY9KEh551k1LYvmbGFopK39LQBUxS9pS/htpxyZ2F51QMNFYVi3w46
cMziVSQpsgUNmkkEEGgGIW1txdrfks5ebiquU4RWsqMwM8iuIwhPxfE+xJrR8+Jc
Irn0VfV2eTq4Rcy8gM31SobpKRAnWAhyPbBanP6Q4UP2gNYD5TDAntPzVYTFHZSB
QFpAa8c7vN62oNgmnF6B/HOMWQ17+U+JPQoL1qekq7bVJq8W4qrORBsW7PRT+mB6
WMZ7VVvG7LnDEAqNrSHWUbb16VOjYkSlbz/8TpAoOXf7kHlYxbLZYmCFi5cL9GTp
pTY4pedWduA2l66fEqyZMbinU546/G4fspqO0rtRlKvPXjXV7FLsNl2fUuUU0zdu
jM/yOYYC/fNEx1k0muGh5Y/LlKNUOQc+D6cgrgtI90kzmjypBokj1p0RSTBd5eSv
EVaw4yguC/1eqsNGRPJkoxzNdd1snfNhpui1NjiuFhlTLC0UzmdZUboGCe2NdZyn
SUnk4S1SZf8vuXX8ck4w4SAKCjn/GQE2jAOR/4pgWrZJV5BgJW7jwybZRt4QSyTI
1QZ+RSOm+CJVagLEVGViDyAyUtjoGNwWDoiiJ21mU6vRQvz08i4jUYTe6X2qEoU0
9gyNC1x5ws3diDwBEsMZ2brSnZMf6n8xlt28aDTJ0lDM9Vu1AHkLa5Oj5DtTaEV2
KAx9/4mOSDb4qq2tsOGn6m6mFSlsIFf8uGN7m0XQVV6IqvmkFWbuLpWEztpU1RlX
7QCWlJTEwXEXEbRIlXnOdO13lKqiu6SSBV+AW4tya4151SNAluCe/m1NlLYzCz0I
MQYTPFZ61s6IlMv+O9GOZiZPp29xZzWz9GiuqJZ/kqwrTfhxi4nWMTn5rBMofeCv
tV3p5AOi5bfWQv8bd+ZmiNByKvMNLm/pBPkydATH4CcK5zCDyNbleeRso8zKhR29
7EMHgvxkFnCgIR3Ay09dYKE6VCJ5V4ieZ1wYtfb7tVFD8DsOgTFdjLfy3sg83hF6
iB6DzDtw41uBt3yoMwV+mqH4oFoHppznhzQwilQD2WUAQId0COWQOpDkzZw26wQs
kfk9RZNkbWCfg67IT9yD2nRekj4MIpF0CFfbQMGzx456+cUYTejiXuOaES+jvBfZ
5uGF7V2BQeT8gomnRTpViCStVgRniZOTuSIAiRI2qryIECjIdmJdfI2oVlXDWpSE
GsgBQNOm3Wu+jKdTRT3DeDZ73IwP/ejVlRbWPiUPrGz3gvHfnX2JRqEZFDF0YdS/
3iv2lPP/Iv35TDKV6fEMIlYTc9Msz8q39/q0+WKLQ38kBbaiEsO+kX/OlbTgQ2B9
r0LQn2dIOsHEKse7XU7T6SwHE0yejvmaQndOhIt5exNuKveNfVzQPu1ZJYrqcrHk
zIvXu0lk+IAi+e8q/ZvRrc8fDFH4RPBoFdLA6RwnXe2Zk2p4ICCGO5ezvoM2aNL/
dbRnJUX9hEpbyMKowMl/To7msgW2PH57m0I1cS7CIcAmIYDcpHnvADHU2+IXS9su
O9xUxm2HYT0nYa6eTpDm1jJ2v3Nyokg97PTujzhp5r+Cad4wwbFLQHAGSZq9sbkE
l40bIFxQ/9MX6DsB/XZ2sZFnkxlWKSfZVn7jzK1UYJWkDZSU0fTV+rCetvf6c4nr
YGa8Lb01lsw8+InK82h8biXW/rRJannVndrjz8Zd8WAg6C66DyhyEONjU7ZUW3FS
urmznUlhZgRE41zx/FH1eY0eBjZZxWm6L0Lo+0CIcgtzd2hjnirIDZG1EsLEOdkF
Y1qB/77eYyzZFXM84sU4evpK4el5OjUmwkoyiFJO2LMwMpekOvu44Nr9gfeAtQFT
dLUWmevHkA+N3zearN9NC4WT7S0RwEsdcZn7g97fGU66HSHDrGUuLeTReNMMaqZ3
P5w+W2SwwidfN02JN65nfbTQrJKhJjvC5PksTIC4t7NHic2a03lV057VBRkdcV5q
F6gFtER6Zs0aRxia4boEf6gUm4FNcV9LgK4cDCnV5PFUWyZpaD0Fy0qz9cU8j576
hDUVuRnkRQDAwMGTU57WhbX87rmTCYE/B6ocUnyO2a3OxBW09DS8P5dLmiy5sIEu
TDR44Nn0KHcgAIdtDI/ngjSUobnf5MWgbRL7n/L6yJ/epQhwMPMrwLBe1wTH3PCX
hXrvoXs6ycK/qGrCLUOYKgvPyIPe6ffteON6+/irBrA8QjMPecRK5yuisbNFBglN
4bzurFIY7MTEHo/v85SlrXM5pG9QO5S494RjTFGCOfrOX4PyBvfJKG8HvGw9lvga
RrIogb4Asc7B/6fQ+2OZx7gm0TqLLl/cX7S+Laeg8gdvaj55lKqUIEIJq/6VDk2/
5XSGCJdD820Uo6jL1qs45w6SVp9cnfCSkOqXrCQG+zFKYVc0DBsATLSNlMYRnx2J
JoGwSSDuaudAC9czn1iszkohDR8dKM5P1YIs1faTOGaM22dF1S13iHKwCGPfI+s0
OqLDXp1MXbxKjCLpMYFYGiOxW7IIETXmJmPHw6mNMwZsmZG9cgN41igJ0p5Y4hww
LoPPxjWjEgHoChaG7lAv94ffmPgiWxc3uwoDIgOrxvd99s8HbOpU0zfIwsknxGk7
U7c/nDPQE140M8YqbQ9aNAREMipQdJh47GSn2VTSWmsTuVqFuuxfLqtJk2iB/IfR
r0st70KnPkuDfI8azO/FkamnMRoKwRgewEE4GqC0p9zuI0yD9cRUb02WmiQw8otZ
+T2193hmFgoVhqFVTw19HbRLkpNjXEw2GEZMNElbKcehzV8kwSdmm20NzjW0FF8B
`pragma protect end_protected
