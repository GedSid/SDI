// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:38 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
O3Clx1Cbgg7QdYesooi6HesltKD7+q34hEe1KiaywH9Yb1lBSS+S4qEwNZ4e6a9Q
5OEfID2bqiznNV+/u79qYTRUauEijekbgJYQhEH1YUJxE3YCwe/qKeQz7bneiHMP
yxpWQaRPAudKESW16rIDYXixZZ8QVnUt/EMJvMLBJT0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28032)
uMStkPolKWNhP1LQ6Vc8MFYor7mpjHQBEgO6e7beiME9E7AN1YQXmrhMaMLuBJQ4
qKGfGZCw2XM/Vg0bkEiflNxwbY8/kFRrVtbfbMKw0LutngEwtNz4nhY49BIF5b45
arLTAIyNtNLq/WXGR3RYNwWRxnizpZSd4FmwSt3d7RFNieJpgzutvgc0Y4hU7jht
LNw+jO3iEOAWhM+NGuB4kualtqulQmyMp7WL3AdxJc1nyxXD+6wqHYdS8IYmMYCx
rl2g5NuuGeBfsmlaKjgOLqwCHtnKTYQdYBn7su6OPVfGenQXQmquyxg2E+O4bfNG
qFV9HT7XYasprnI8NuR2PfijbU7u3MsKbw9gZgg5GL8MD+qcL5N6a7phNYf55i4x
nrruVuYBKDnpb+9Gp/ALPURi3KH8PRZDCnBDe8F9iCew1PSUe+eU4oOdXckUcxB3
EGmCn5rmFTeMnuPJrMtrxRHRPEpHR5+TXAqzO/kDWlX3Vk7J2FVpTQeQoFxQ7Bsj
72jXM2AsjsUc3TipMhJASDq27DpD8d2OwpqhKdwbYxJoJIUjm3sxCrixKkrncApy
pvQRIZqklw3ITB4D2clWxyKUaC9Hyb4PSkfJnYJ5JG9UYbwy0hycsGr+MHbOopAS
97ZVlXCbzExGgjPAXQS0X5LXXFDOEhni9edSgm/Rc+sDNiDnxlnlCnSG+IJ2IqvE
ey3RqXMmVUy7957PEXfpxjk7BsUgrPKvhMKK308TiEh7LS11ERa3QqGZ2O+uwTTW
LNJni7VXXxu/hlt6dRi7w6FEhySoWZU+cfJaojHUonYLgdA4n+cuwVrv7mO5q0O/
kw5Q7OcbI/gCKdD5cSSikBQ8QOrya42HB+zdxWC34s4YQ8X4WVtKlu7sTTCgZGfv
+hXbSwk9uGPCzbHk81he1Yhzj44kvwozOD6SV3YYAEJngy7kv0l7ott6+EdARVtE
tPjcPKxIIAKhF++1Y7zWaYNUIMeblz8l9WLyyZK9F6fu8TTHXnWm5N+e/0Wwib30
SM5MqNsueRNr1L2GSEQrjXpstG+cdBfLm9MIC9tIaLhKB4y0Reui+IAgHmUHA8CP
2wZIBp2ezGrxjJgN2DPzZ/7yp0ehCnXmNVn0cG0u+6Ki1gLND9tyUAms1ChfiC1J
vOAFBTjIXYFq3/oXHtNN+xpDJf7piBcAeq5FXTEzP+YLEnavAJajQVnc5Y5EeaiC
tSorLNQYN0lYBQDgEdlq2mKIkuzjHV58xkPxu5i5ieAHYdUg3rRYFyzzVZUlY+qA
nDj5Sk+v9wszdXwUQ4ghibRk3OeeeWA54+2PL62YHrT0SSXWeXfeKD5BilUZkji/
+pYe2UyrFWE6+d1AjhI7Xla5wI72pVRDXVewRqcYFAO2s73FwcPAvdsbL5aF1e+h
jFrQ6afcIpmbptIscY+NYHOjFj27PwOx7Z0GcEgTxUh933bST2LahrPrxdx9Eewm
pgISFJwxqGltivq4AbZNrxh5Ug/22aOHn7sB7Qkde5ij7YxtsGQ716aq8s1b//ax
HexqpyI5TUoIppHcivfeVa4oUE1pdqVkURKx5sSUVbQji6Ym61uBoAHEZUY2Sf8S
A1UNG78QV+VBQT7oUVM0tnIw1qLClmRcGNGGn4VitJw5WPKWFFLwtt5KmL2YEnNE
lYbVePkHDFyfScOuCaKfMZ7sMtnP+i0feODcXBf7zTdQ1i+pU0Y0kG3JPji/iKO1
6kEtRaB0Xv9NPm2tB8X1Pk2mPrNj8E28GiDvgdlCJVMqBLfsgKSb8xspbMmXIBBM
hruz0DMIV+PSe+aCO2a3XjqreXxdQal4r4DVdG28F4UkPljC8lIOOGacCviKnaQ9
oji3so7sLmeLLVLXYpur0qrtq3deNUmNJsoiP5wR0gzZYjmaOM393A1nmzcayshT
UttygQ/ZsWY1r8+pTZdQOlXY94KhCRD3y6rTzEiGvG9jc87gNPSmnBSot193/iwL
wCLH6KS2AW4GCSeXuamDT2yQvWF6iH8c3K5Mti0QEw3QB5Ldrfyl0HsMINPWRfVY
clZ+KYbDniJP2yRKWvTXaKYJlk1QPC6RYU5TipSnsXQv9I3FFeF/vWszXgUFZqJC
i/zkCoBtqkdEL8mq+j3Q3oVE5EwFDTRMWbj3/rhnNEKLdlmrwaw5cCM3mgd0mnz2
t2s667wWIWvNIUXSUR95HkiXTjtucjJwGyW//WMc7iiuwcLCnYRdeOs5ShjIv3qC
P5vrvdHkP81xLswWLz0HqSs65tkxaDjS0Vle46f0/s/27VcRKqSvDQ9AXe+6BitE
AZ9Kk58vifRrIu9K73tFJwE7szTWnRrZIEZeqdeT2eQC8uL7nEWDI0EPXi70wA9f
YT/1YyMp0QcqK++6TnG/7N4enIuAYZ5ikyt2sbp+T/be+zdipcq5hd0n9fmoIIUc
RYcI4bQBsxLBIgO1JFw+RDFD3xjliYrBaj/5ek+umSk+9/nPL96rffLu7PMedBl0
7q/1M2mmrUG42yq8rssgq0o9sskwNIM/tfL8CtGeuYElxlPDe1dqZTtip8syg/gm
P8btU0LTyBHnzaxvsJCI8bOtMkImag0D34I096NVt1XRb/BTSygsWxBJPCcXadAn
iHmKGwJHu8ZSI66hSr8Ddrt82gRyY5m1iXCTFo2NxKDDeFGwWPgBK5W938BiYT6s
4pzA5G6DCz8ikR38NPROUbjcX5o5swftfAzvDTDDxUzlgPckkLr5oEERyn8SW5YW
z4C74uFled0l7ETKlPYJJrEKTbj8NZyM8njfoKhvaG+aF0oW80Cgxz4ug3IeqEKC
yh2PQW0998n+G0wCIXL7eqfqP5VtImganb8EqkvMcAXtaaO8o1B/L45yWImouK3W
vsG3k6sHzzqeRHb1Y8+nMUhTK+KT54CE43SQJy7CsBzv/PWoVLlMi7aQkf9WXD5L
I4ocG0KTLagLAmTvGQ+9rro+E1GxRjI94XCUfcPQm+JvtpP4Hzo/k6s/zZz67w7D
B7a7qkZhaKkb2yGq7Ne7M8v0TyqTOWiiJvqBosB7KR7qgshEpaWfOc4xNQz8SJ4r
eVASnB4fHwu0GEFxFQC3dVunuy/SZDIZVEbA7212ibl/AYk9ggqmofSocfbfDEtR
ax6zvipmDuTNqgnqNuf4X+B5Ztu6uyDcwWFNxN83sfrKaerOux9S61tzSCO/sX3i
CvQOObu5guqzN2++g4Ge3XrHlThj5E2kG85HGkDvt3Z+6O4I/CeT4XOuP90hNXT5
oR76/pgmts5oFTIHB++VWyf0eSbDHI4BoviTLbpdvSAIhRVbIC8+JVE/0RVZf086
5YsNows8f66NN0jPqXA1s6i5CpmnDeNxDbKH0L/u/gyFntLzoNEcTzG2JVes22kA
noDfKI6hneB1UHEzKGl1pIbtLRCYPkeoQPaA5tColduQiju0acSKlSSL3rrQjJf/
6UsN+OaN9+pSBBjd5RgXr9DIE6iP55blhvao39+m8liusdg6NNyi9Q5SlS3EPYkk
Xj/A4NlgHsAD8xza3g638SPO2H5AwMqXaUQKd6Hxre232OBnw2Q7fQBoRou74NsD
ZU61YnpOEQvyHUR0s16TmdjjiFzZ+avK6LfkdfIGLfgF7jR+Ny5cOy5zUyWeG0bD
KiiNwKFyG4/odD32kaT2lR0qLb/DzwoxC+E3IyPLVT474F3TiWSNHTLh2RPLUaFm
7ukYqYGMHkZ93h1wCRDjnR1yOhwzit1SuWTHVR10EZuqbtBeAy2PP7LqfPn3sBGJ
gLcviMnsj+owpt0hCltiWDxKdR4gtgd6xvZpkvLStVGr75zSOFPvbRT3l47cqO93
PDPK+uidFul/F1D5F5azghJSLNpczHSOujdJgZfinT6gtrAU0Ibf6fUV22zL3RYC
H7sEerd6j2kGxoIhI8JftGMo+/+woIJDrDx7hDegpKNvXArfGuND4myeRhPBqJ0Y
w7oIbdNUdvgxV8eooxP+aL0iG87jAZTNPxPugH0e9nMvQvg7BDdeg2iz4avr/KP5
zGXJe3BVOdFzptITWKwn1Jzu4kUma9MwZvJnqRHSs2C7u3QV1Bq/8P5jVOq12WWi
/1czVynOgePEZUWv4KJTJhkmadXGw4raBpAQAIMD2mTij7qLznbBSMXM+GubbW85
ZZuVMuTAst6ZubvX/5f3VPkbxWI6vZu5jBZBJ+3dZqz8FtKWLiW/B0Vb01ucEuei
oSCjXdw5ken0oBafatIujgsW2cfVl5XFr8rQxX3autXJQyRMhp3zrqQb6A4Oxerw
nY+acL/+ZGshSNALBfuKPtTqMvn1HwFczsGBHqXg0G3cWFxVX7hDITHdZmZOUavA
0QgqeKo27wqBYCdtCGLx5GX6EOD+Bf1wt/vRO2qiojTDqGMeb5p/bVk8ExKegNLa
Kh0YDLVJ2GQnJ7JKr/6fEJsDkr6kGva32sxQzRts2eVkZfDC0XbPyLA6vRkBkJv+
dnKOnIiVCfAXeMsblsQ4GuG0MgnyxRbwNWCoXbCrYmURVf6Z9VtULfyi+6gB2VTl
5j6hK7VaN/sST0i9opWFoZwfYbLFzUmnJMPyOFIEa1X2kxsVSiQpM0j1tnHkJEEc
gYDU9TaQZCGfBNkDIcBGzqEDbJs8uzezyPoLUUfFiTS/BonvIpIIWV41QFX55LZG
d7yJqbL0FzyEd+2Pg6fqNEolqG/27erkC0FxD73Kh5NXJnxGMh/kro2dq8Oi76t2
RrXbE7qVuvHA6D0uTaAMKT19vVPOOoMhG3oGI8ovyrrgcRAFjctPTWfX7R08MP7B
p7M9Y748V5VWiAK4buGvuNdxAek3pato5Tazu4CiMSxRHoz0Zr+RIs5PZ6qOT6f8
ipbwnb8ucyWWXoK7fQYBAs8tDsGV4d2qLifQ8faAmlK+4BoIDZVwgz5SP6woGYNl
A4Xc5Ix5mbnxcQ3Hc4yk73a3rnPTPLrLi2iurgAnrywzGQbq+g5E+qUgIaOLPCWZ
aDvebahwUWTEAm4Z3TD8V/0bOZ0jJIxB0VuDbNGohQOsb+TOltC1V5Cu5jBB/j26
19PCiYbW3vh6AKBBcbVDrQyJHsWWq8A1H3z4SF1BIIyiCbXkMls6FZoCkTh/oQfl
BAy6fviD4zELwKcdQyhvMTA6aompb6JwAZZxSNQoyBZZZWnJ0T1Zqvek+QxUxU14
5VtfzSQSoQ3fcq/3wzSQaJv9M4R5naSmmTzrEuWhHgKZ/YFg+inTLseAFhObTyOB
rv/8UIU8J9WZ27rMbu20CxgGclXYNyQFiwVFng66Z2AM/nxS4AEH8+zX42Z+htaJ
d8/PcCs8uMdo/VX17noWsbdZfDRUV0Oi2nJskwF3YkKCAEL1hd/oKQDxrOtgCUEl
1ta8oBhKpdoK4sm+JOVqnFdbHekl+6es79WzujoZaBs3lusYQS4QbLU29CwDXqfk
LbcCSZFm4p7TfWNHTiTzRgLJGipRmg5NHTgmZq9Z7UB0v6PNCYQv4vn1pzKseKsm
mcVFgsyRVeinwYhEmT5NHciFw8rivrRiQha+SQQTrUOXsGI6s7hX+CLf0Iv9+Z4z
QNfjsogF6dFYAZ9jpOt1FfdwuJiZm0CO594kXt+ZqUBCtEsJb1S/4Uq9OytDR29Z
75koN2yOJEJDq3LlZJpb7rUjEhHxLqiF5liP21H21Ni+yKOk471hXBmzm0NqrOQE
8dTc+uiHGBQJjbyePn/8UUNzgo+9/Tgsj16R9+FhJzbgrj7+64baORUPza384KbN
x58+LHmtF0rcXwSgLLKpfoOIqvzTt2BB4TfF47ILRvff882hs3KbO8vs4s6A2AWZ
LwO7vPmvdCuERaBMHZB3wFfp0KL3NtVyxTwrhU7+NPAGp2kBGXfAzEGcx9mvLHWa
kTP4g17gDXGP+2vpGqyHwP9+g5V3+UvWbItXZ7KPMo/fwYJ3Pr7fHk4ooVenU6NZ
aqa4SHBXJNVtBD5c/qRfEQFkoiCCEZnoCzi/2DzQQyxbAgp7Lm8GmdQpUzOkvPjy
sFiD6B+p65j8NhpoZn4Vx1WMHgGZ6J8EcQTCbsV263p84Sf0AREs7gqijHjN/LBr
bnv061eh3XAdJ4pddKP4fzIsOGRar1NNCStGvbQJZnkneFUFbqSWG7mD3kgBrWI/
m8koGRG7Aq2oGvm8CqIxoOEQJqtOkkjylA+qHi42Gt40VcVzSoz4KyybAXgFacxS
LyWzqYbzzWcUwDB42huZRjLF6qZdzVKPCML0YUSvRJTLNiKdpuoaYHYwBdBMV23W
aB7nIA8PqyG5BjIJCf9EPULEdySUGXKxwtgFST0d+cnQ25h3GCB6kK+Xg9lpySya
iDCDlB/XcP2H9SkFzKsc4X8hOIrEGPccWxkjYdJHhZiQHxS5iyYLdq56r5Z9B8JD
2Xse324bYSLE3n/nGt/mjsXdViPxONmdYD+a7Puf5mlrr1nQOhSQWQCjRBD24Cpz
vtamsyvdS6ib8H48fRsCSzcLBB5yF8P4T/JntxeBpjVcBlgbgZZymP/8Yk8uhLa9
c6U85hHC2yucPV9CSY46JaWDKtQzcOt1VYPgyi6HRv6m3hsC+xvXmwV2TSMb9B6R
/PE7Z1AnoqOOVR++up46OKVs0MnYblGBiXNgsuAA5u8quSSsupcCbg8sfOIPy6Sk
zqBJGZSww6C8KdQeG+QGBCGqwn4EYl+fmZokTpnfcfDlTHffxV0UAx27JLefFmok
4Trn/RKP5y7nHP2iu3BK10hVW1Hi6KJ1LbCWWNG0qD/BTGa2XsXsPIeRw0ufWXvw
OoDtQywq+Vq+k4aqPryu4TdvZuAw15p8VRozKAeeHc2y5+waq4hLmwlGq6piGNP1
gB/tjb3ze7A1ZqTL/BaNPbpf8I2HahwlC2kNiPlYYXPRUVE+5O3jOjInqnosZ7BG
XFSNgNfD10KDzrF1qcu6pjhEltVdJpYcohuh33yjw4Pc7SJ6DTzGHBpv7AZt+vtC
S2ycNDUfI71WHSdt3zU7Us1X9UA4oVo6oevAUIo4+2EMaorgISMxC7OYnWozyzHT
nZJkCWpBtvVLBSJ2yihlVFXCKN7khsNN2YuKCvyaRQZj7nfWmeMo83UnS7Z5B9OB
f1uOBwyaLH1ioj6vqhRvBdMJpqexbnbIzzB6nGeqJij2rjWt54oUHf1Z5/HyNTPW
go9N+UyruLeyp7xgJkbYnuqrCxl8RAviRqVfXcP3wuMUASrFYcxXHO5g9uv1h4E7
oabuJHvthEP/8SmacWzmQthlE8Pf5nbt51fQ7Jcs5ubV5hnFSGk1c9LJ1Nnu8LFi
2htqfBVYj5k6lzdgX6MpsPPkdlA4QW2/cx1ikiK1+k4FliYRBMq/lRRqzLPOIhhz
KgN/A1DLXT11huDdCdLPc0M/Tb0bgw3CYvzcjzTzAWZ2+DG20GtKJHqrDa46JI0e
mlftpjX+UbNLBJ4m0eU2Cc8yk3ZDF9NxRok6zQDixe38L8gLLn4B4IhIwdArxlKJ
7if/1CEciJrtd/AuWWCCCwIOlETyfn8sLVWtMk22zjQ5g46Je1C5kg11siX/8Eca
Q1hMx2XZTP9L3lgP2Ga4PfusyW/ItmK+t7Jc15Tj1/Mh+Tb+VN+yK7wHdBZ3vDdw
HAVYg9bvBdhkvDgC0eC+tXted78qsNTkFWgwhRJBtFfbdIqKZJH8RwiKuWts2n16
g+ZdfDlhxUyB3wpBVcfsO/yJPK3L8HgPdhku+OC5gpX9lX5mX0U0L0a22MYYFKBS
cO9cdl3dbh+LtZZjm0eGg5ETF8g3dsWCVq4t6R4sK9ZVS/U7EP9OuyvysfHr7jdf
f6gonFTIJmCBAy4UYE1VZdQcTn9TJ93lx7VbFLXBAGQvy36vW6TIBjmbik86iS2r
llz075sktSia0e7Xj81HIDJO0bca42hYPCLGaEomy+K/SxZm4J3OYHG822wZrzYn
NE6SqDpMvJNUpjs1dnH1qyBEfqRGyPSm/i594drm42U2swr7NmOQWCQdD1R4o7Ob
UAdNpOXrfBCkH8ILFGWmuc+jJ2Z0Pj+PVhl28xyLnjf/jk92dI/tiw5hjtKS65n+
hUa2RgXmBtH5eaWVC5ep3iwTLvfbisBMpsuKghE1y7NS7hBy4YxwliqDBtgBM76N
tUYV6Vp0FEBdTMdxevIR+NZOlQovxAdfAixGqz14Mom6jHSFTfs5H3i7DICAPjnj
efzPLbuH3PSMtgUCLyKVTWFaTHifS+bTjmcBdDDeSfqgZ58ujqBWffeXwZ9Ic4VR
3wvLTPQEO8QiOIZW0lmPc/U7xfFJF85D2aBtYJ8fW+WzbaKKDE7/08R7sOeej/Qo
DOEgfJOPmrcaG+PvpbyCnsCHgbT9QgpoBXqnW8BWHLTpa+8EtAMZl5gIhJQwUelN
rqoQmAH46etXDcAxDEKpviRIz739nikkFcX9iuqhQT8MIJi8+04OqFKfn/4ay9Cf
fTja8V8b7/maB7fb9dCyTKh327mVbWTipi4K6PRlV6pghLVILzEQMZ6IiAGflkdy
zvpaB15hhcYy9ranvPFV3sfQJJULJ96Q+Z8BdzVA25yZxZynIULzV2KV0CeW5V0l
+qCAZ480n8lLBw2Wsq1g8J5SAvygwnGw2q3Mw/PEVYDliG6LT6Wun9ARvGBh9OZ7
/sk9QHXwvvC0fKpSxs5WKFDn66YopwdolxjpAbBMzgy+Z0Q4RzYU73A/XOgg8itX
NsBxTzxaJBs/nX6jkjk6owcj64G9YB7z/OmskiimPm8HtsobDYpIWTS+fzaSGc3q
D91RJJt4BLPsJ3ha2+ttG7dmaE4+w9IAP1BAGn+L4vhSMTJhWNpakxRAKsASoan/
7pYhgRjwTx7wLYGNw+Z8ByGld8E0PJtuimB7J8+x5Ki8I0FukTbKNYMulupmgryh
a0yZmzwd/g1m8+sqIxBcZkoZcSVaQbE360Tp8Gg7hz/luqrAxZVs8Oqb/io6C2Vf
G7Q41g6qC25ZzUigENtWYkU2hSZVFRAzRcB86EMzWuZXU3J97MP4OfhoIEg5tULa
JvrRDViKdHfmxqiWSuOzbtxH2Rfy5tyDj/EC9pMiDQpNdD3oa16226YLTUQufN8v
UJokOHAcfpuUolhCEp+hkJzZl5133L53M37o6o0jHrlraihjoVZxM+QhjIS+odkO
NBt1EKpLGAdIA5rfhJy5b7Gmx6XURJu3BuI/WibsrSzKW/tSldajPBjT7H/t+qkt
5Gn6pV5/lOyag5/CBsK60mJr6PsTnlUnhRf3U/eBcNjv7lgucAGa8WA3TzSy9grz
FshPQqp72MNnIHAU/BjOqRDgMTNKKQ55vKBxtJQT3NxZok0VlYTX13JYE2iLdh3s
uoEb5/jYyjHCBO4sM4DrSZpQxSHIGvvBJJ+LxJB4NHtOBjqXCSRAHr5/g1w2/cDM
g6VwAnnnwkePDtkE1OegA+yOHG+a0zF79n2YJsxSkvVOBQCxhnFiD3AomVA1U0cj
upzwIaT7a/kCOwilgAeqnSaK5TjIePrqj/hJbIIgnt3cmnt8H+poMnuxwVwoII/s
YHweRs211q/BOfk6XV8pcm8Z2c3ELluXnQd/e3k/o+8uuhW9sXCGkmZOR+8hNL2O
J5xR5FOxVBSIFKP1Xy4Z2YidqMsHykymA3q3Jw4FTt6Ar2bBdFz5XmI5nILY38op
1mYHtkRnOOnwRtVQ2l7qW9fXMpBpK3JLeviFP+niWx9PuLR4OmbBDqcmgiwRi5hq
aifK1XI23z6JzMKr1HAxyi2x7hvqWrXDKtuAx3/FReUL1I1tEwYreLCnqU/c2Yew
BofdnnJ7gp8NOKVy5tQOMxfXnWptNBEBMdB+657/IC1dwJ7mXc7mDPYAZ1ZkDYG3
EVaAwLSlhSroHPOQsZFhw/o0MLkLMC3+QMoMH4CXWesibBrG6gmmp2Ztf/aGYZv/
vfREt1FBuZbjxpJJ8T76Idm4CRQxf1NhLDKntTmJamJKDs58J2t7aWO9mF6aFZsq
sXovCqGXBl66MF2QWTbpR7uytZ1gV1Hi2OqaMgyIu4OFbkzW6uQakMfWDK3U9xFd
juowJaNCwtK7ypCU9vVOs8YxIdCb0CXjfSvxWWq+HX0e7wdaikkDZ+oLt77893en
KLhh2xAYMY2Kaj0ChDqjo/cETnJ2aUAW54AldpzWCodCWrAhn1a32kuRJX5s45+7
9QNaRM6PF/EqzZp+qiIMDXMy1zoQHDPVZb396tjbZXx+611O2awvh232ypwawAf9
MVfNAprhW5kgl2/LVCFGbByAfc+SpHcFAlPPz1C24vsIUNKQq7N+AXLznhhDpTcW
2LXpYjVrWKf83f8Od1AUe8JBjuG1boKg7JcznAyDVuc7jfeHbwBSRqgoReFhQZ8g
OdmqJuhgTv/Jp2+bJi9tzyZdtRBddUNcm0b8pAKVgdJTtLrEdTy8MQXfuLqIT1uF
b7PMnsHTdVkh1k1JrnmlvLNnFJwItEJXQZYVD5TJ4UvxS1ThhVZzg3jvquyMvPYk
i6GwV1+tqN+YfSHhKDSifI7S0+Tf50YFuf7UVhgPua4iqRKBMiAcLMkNcvdw76gG
hU/IBA6tGOpsZNmFV/olct1U9MpvLLdUtg9KUVD3uy0mYWNxkk8qP84IAIig5G/O
Qx48F1SrWXPYdqOjgx65a4B9OWAABLo5SPn+4ro8U7tjpgYqOAXxVXaqP8mhEkEv
GH2SlamxfxXpl9eHMw3joapE+Tk14C1BFqzHFpGXUScvNi3rZm96n9z368OZuWeU
lPybQ7YeI0sNW6/2DPRA55IWxaNHMv486CmEDvMyr7oxT2+KDUELop4j5wyCQKDK
ZgG9ej75QQ97USCiaz8CQ2Oiuw3m8NjglceHDyPfeq7Mn019BWnBGe68YzYcvYmz
ZDejcpJD1CPPfnMB7CoqW6bN4BWDZ24GpU5HiP+dpjtzcIui2Qw4Gcf+PYKUcPDj
6Xs01dtOEzwQBTge5DlRmLIeClW2yrLYtWxKiTK/WSo2qyX7DsIt68XbrjWPh3y2
aFyPr1EfPYJtggxh6dhM6xXQjIM126V5blHAwlqCzbPnnqiJDRCX+WqDtRgc8KVD
S7NntJYC0ueoyNRkmuVwy2VF5TlGnU/gsEzFwSW9igmis4+hme8Zmx6ccGivbEBi
uFpzYA7cUFHhICIEVwKIj1DFxvPzD1ZG3Ffzsjo+bYHtqaOFK7MPxB97UedjuiWL
tvzuOGVSFIWa5/mJyiCJ9jHXinrDJ99sUVpSZ/G93VJElyfEGsG/0oMf2nn7lpxA
HItKChG4V1oWx6BI/1WddyhSeceoqFWiA85T16JCfeQIq3TbIKbJG/WA9KArZW8J
XZc1L3e+urD/KWCzHZw4Jy1XeasvMkWscrAGSQLdelWeUfjgosQG6GPsMDKo13dq
tHC3Fl8PSKk+v2OPR+P1UFxsG07oed1t0PCK76bbOGtyLgjJMhy9C/e2aRV7j6Fz
2NBkoXw9SYqjCUEX5ow2XRUCNLXkNQ0deMD3wHfCMafVn1baqSb6BKMdfxEnhjdR
5bHC3Ynt/ZkpClP8f2AiVhzGRdjYiitr7WrXzsM4R8W8igP9tc35OhX4oXGtLHll
bFIc6VN/0RMnbF5WWUdU+YJ5rqObewpQh0owNQ0AhkcwJbvtJ85pX4xsjeCZ/aER
+iM4jkPNBY3jo+QJ2Mj3KnW6ieR1gmEZL8f7v8vuy6UTqhuS9W05Ljqj9sKQ9bcG
pKyRqHwzWRSbrYy1EBus6yqsW+mNWNpUPoGxdXIsu/DpTm6bluT/TIXQJDbHZ1nN
x0BJ8e5agooQdlwQuumh+Em5BNr2Lvk+3X+Ifp4SpRLFyFPIB3rfTWlOTh1kkFdW
IcPI1T9yMp1XM6CHLRId+9t/akYHTtuYbAN54oMMNqk+MB3tS7P4nRPRCCMZ+wQW
RUSUBOMo5nHKuqLxmpb1aaxtLZpByE5bXf3W0urQWDsh2xYUL8bli6Vcq5WNGYDp
HJnYe+EuQUFAN+EbvUqXxRNkhE7zTa+N0OKMlGV4PXZEiGQFE7mrtNWptWHjYSL8
Ri6LAaJcIlWvMk7duKTE9WGE0RnTZTy6gd9BGx8pR2GTNenSdX4sQu0+haRsR+mT
VqMkSqn4i5HStZD3vGug3nP9d85ykRKGvfyBYv+W+Jkop59H97OAADskgATRUBm0
Smb7QVR/0dLMaSswG5tqJfxkMlKaUeNFrQ5fflky3OhU4mV6WdlUdrFu5GRNxPpg
HEPBaivr/FLSuJNhA2Vfawjr1tslKwaJa/F0JoIAy5NG+H4P83LwAb6DPr8iBnMD
z4ESMgOAcM6t23t565GkBakGHk8WvvKet5mGMtn+CDIoHpmBZXzJjzHKfzYbT8qf
+u1W+kuw0D6yPOMRpBQ1hSfMXX5QQV5umo+a21CAkys9G9XpszJyUln4bXkogibv
A6Ci3EuVoVJN0h+55ua5kEq3iKPY1NBOrx69fsn0lYEIQrHvDjVxtfPt2sXF72/n
CSUyeC3U03NCEvHYCuqhS+fwsilyj9OCP1VbI5OmQI4jJRZ1G8FHCXhRTce/oFFe
/SrHVSRzcRVhR3GaJoA9n3nfnYr99ryDLdA7U+N8xxw8sd4jVrfIyPZeVt3rd+/T
KSZLhVn+NDB8UBg/UYQRJgDN1yaiotYoiN99/tQmr/YEy6DGjy9eQczr/c2T3yth
AVlc6n1P7poWourh/QPkfXc/UiIV+czl1q++svVJZIqmGPV/G2yK3jD2XaTxWtLi
on5ssuUg1Ip0ulONX5Q11NIINBqeeQJ5MummDV9MdpqWdURv/0o5vVapEHhGhY/m
v6dlnmq1drs/yGc3uk0GbmiidIERH/ELC2u4qGBVO34ZO6kJIaagpgkVi4K7Npv/
sFajd9dJuHUyocsAQMjOafUuW2t0+sZ619Pm94Zro+JPSrOPRYLnQtlcCVzvHsiB
0lieaCsaQahjFvU9ilCzM8nGwxXHO5lqG7RzlzuqAHLl/ekHXCtC8M+IJ42T7QgU
Tup9aT/pERQUEtNSIvYcTNnNgNpudPvm4lHBfdgCqmZkcPIzhl1rGmQO5OC1sKbD
TvFsITFZbD2euroqMGiKw/rv89+J+FF54EYtC73e4qDFBuGkf2twVCv0HJao2tSF
2iu/1QJC5ZYTSoM1TUrL+8qHcSq5GdNdXlpmuEHuC746XmmjESi31ZAMt7UfFt7g
Lv5Jg8kTXDFRL6oWFqrDlKDgmv0ohmdTxUsF8kpwuAm1r+NrQQRuCk7j/3ApIjNg
94QvhVQvpC/ZxQZY5Mwbc1bqYmiNf5HI/Wq+1pPvvzIvGPtljcpA2doFTk8SfTWQ
xwgcxZQzrdrSVzhcacxOlhR/xsqSWoCBQVNwDVHY0UcO8scaxtZT4m9D7Cyr2EcN
Wiof927UUjp5fRzvtO16EUuTlITkfD7ITEcokVfChLrc+p7gcJ7pic1QYa2PrtMJ
CL7bl+NEbsBB/QEjtmz163p3uSGDJXzBqYSQvQFGSys/8ETtwkc8XYClunZgYqwC
IuOSfZeajF6XXjwVOZWysU2N1UHPRSGrlInfdo7uJDc6VBcYgEhGE2YrZisq5VTk
2LklA6EiQdjCAL59VTMp4YBdBSP7psv0OJhCfnQp4vkcwCCyHrpXQ1OC3ObPzrgg
QZFEXT4S2ug8yAPMbDSD4QS5FPtsh02ATI2kxQG8eDv4YKCX3f+rD2//GG0T5mra
HgF2HEQ/SA5n77VvWjQc9i+9VbFO+gQNUoPw604sRg+YBA+iD9EKtfx/KCrD8ko4
uLEx5yXPd58F/ZjwKaM/LXs78ch9t7KLs1BCVZqHQubuHbFjqB63078XSuj6Nrti
pwCpfLittaCMq/hh/RPBTWJPszfxyenMr1TuIPIahoowIuRVC4Pozt4Ge8b0DiI7
z8iRPrv6oi2X340SIlYnEc6okr6+gH5OIFJ5VL+TAaM+nP9wfiKcP3QjisGLfIBx
OWXECaPQAqNqfjhRCmLhdlY56jPbqHeIa7xToc6S1KyEYOWfvcxVfVweWAUutCb+
o74mg6u4sSrSjBM+mGTUEHa8razgl6TwqAVdC0z6ajCcYlxLgw9bXfl0jVt3d0Ze
97mLwItDW++MY04n8ZRopD2H9BiRZhMV4OYBKwZ/YihtsZYy7+T/rozLV9YWYLFs
BiHCrLYULE89B/KGkkiYS9hfFISAEt99lHQ4pD/nTl5cx7jhYJEPVJMisiOeAH1E
dexO6dLv3xKtFWi9ofehKjS7F9kOEIpQ9KK/jHtrM4BRMy57f9oCsfTAktZRNiFu
jsmKXg/rk+NmvrdRhlgObDcISnA4U1KGEB3+rN8M8Dh3gI+jFsY2J5DNxwe51feV
oYBzI3FJKrJ22aoEl6IGNVPvPDAynIJdc0uyFJmzM0+MI90uD3FEfuUD2wecOfMB
0Rd13P5R/RhI4aFkRmvGFmhNfIXyG8/hPt3jem38NUdcOtTZ3hJdfcy7MYNoLChL
4VmSaItCBMO2WcQkOmyGqXm3YZa6WanXKhGhU/rTYjXIB12aQEeJE6Fr2z+eFlKA
F0ZT3HSX7Ud+4pZRWHn3cck4Hxi43IPFFzdnfjyF59B9a2F2N9cnAfQ8L0uzlazD
gb345LWSwJVswpDWlyi5TudgmxJau8NY2ijAo3VgnrLObnj05uULL5WBqi5Nq3kw
jKUtGgj7DlKXoCog/HRNkAQiQYW6f+24D3HvTykwnO/Q3URfNNqDErugN6lfrEJa
s6wgNfV6tNdWKo0PNvOliJ/rv1p/arO3EBhzbJC/nNlluIuxdCcszjtPs1tgYiTd
Z3Tb1B3AeL4q2XxyX9t9B3ytGqnpo0ywLE6xAFfK9EpqRHjiJSyY+qfXzbe9aOT9
yogVpyUfvbdiPTtSMkNaYszbeuI/lfUStBsKuMRszsAPotcSKij24sUO4p0TR98w
FGagmQpC354mAGt2uP0wzqv3IUyT3Sbsb9RUGQRMF4rSbOZzMEMw2wixi1KgsHiW
Rjg1QEj98JUS2MeP11fpGn1ngDVDGbKcXq2wIzN8iLdwVf1vi8bwgo9k7vzfP3dZ
6N6c+ltJayhBJHrdOroGUWIAs6BGIvvtSUWpfutnV23E4OM68Kv9K32ZjiP/ml/s
sXxpJgrL/3FNs2HZhwlTF/WvclDh63ccnHbND97zX3PipYNL+9pD5+j3p4KieeOj
wPAdvxKbFMhus+PHFSfFjVeftp5mFldy2mzKS/k1IkIz207GfyGiAqASckZt3n6U
wRyaY9XjcR0ZtTEgtlHDfrpbNWRmvgGh1JQt2cj60k42LXIMLL+8Y2XTxUTlaJU/
seYWi16mItA/P9lmvFBeHG7HnV68m2OTuvF+VQdAHgUwKhfZZPrSToCiBrkN904k
5SdCTF1ZG3THoN6qBg007b4UScElkfxgUhSsMMHZJC5wh7GUa8oxim9wAwv8+hxT
hceCZcz9SfznP/7m56ZNYxoIwsKcJ8b4cbTX4M8cSNHOXmteayiGsVfW2SiSiPh5
WVPVrqY6LfT1UyMAab501EFDC/GheDsJeTO86lNVf043YgDoUDMmVSq3TgsSoT7b
je+sd1sHmTl2MA3FicQ+KB11w4rHLLRWVMJWH0pnlZne5mYOxOjaoj3H6qIt5Y9m
t2Z99yAUljS4VdYVjf5CGnLHri6V2PLM6OFhDu3E4U9L0a9s4Zh0Uvei9VWBImVi
IXMH22dy3mjxRfApF+XSd8jcexYO9gdMiaIdeTfNzF45R05WwsSNdhcpAS7qJSKa
/I0Rad0jTi5emif66uztVk8URDYCNdvMnuWq+MWG88Zo0xbwSEuwj5d0Bsgx0KU8
ygxTaVAl8p/iRL0PxXHh/gi6sgSAU9AYCb9oWBKjW1LOS8LalNiXPONSHSm/6QxC
AqTEGD6ijLeO6zRe8zkCwomSwU6kbZG33XelKzJu9NYkomyguPZ8xZ/xM72U2RX8
CwsHi6c2CWS6T9McaoeVBM+j5w182DMQ9xlP63paC4aR5n/Jjo/rSDGrjqYOYedC
YMZMVntwuvGHS8KCPsBqj46GRG7Df4cb2LW82AcN8jR7fCg6XIqOMlQCeHlwgge/
g/0Z6rEwIxEX00j8Vd47Ews/X5/4GWVBjeePRijVFZd3q6gETV7Nl0t12j9wqa9f
IMdIpCpLlYEjP/UIUk2sm7pUH2ZzpxswFF0isPaLGuqbXmlTCYoSxfBS2r1Sq8Dn
VU3uaAK0mWyza4yy8BUTQH1SqPg2ldpB6btI2xel0ObGfEEQtfktyIQqTGt3+cHe
mBmW5Nl8I5eYnY0fhtjeoFOpLv1HV8kfnIdhPEMycmI6orFimiSz7DE9pd9OgdLx
8yxd+TCOL3zTY2gRAmeFwbcF753hcwZQzWzrm5vZj+WMTgOGIBa+FgQ1r9LJA+Ax
Ykw5V5CJzrFwWyyMPCtBePjGrlb1R2uMETmeO4YoHIeKDLa/PpBYgfXTKhCQN4Ks
ECMLsRPp+d9nAL/kSo+rlHoOFl3jG8GoFMMoSmoHwGUvg++98sInlYxmy8JGcW77
DOwRLXIivys8kX95OVZa9cJS86IqPPAaepytoBh2D3rB6ckJNHagOBaivf0Ybkyk
g5IOht7p1ibBF+u5f1c/7pDP+VJCZVUW4Nt58dfMpYyElIMsih/KdJ/pswKPCAu1
2c6+xJEY9k3P765w5GsPhkws49/ta8qbtbHbBp6qR3ODYx8+yZ237/uN3Fx5JyCz
+N7bYtJn5sx+2GrXQn7NvEg76l5FGbY402D2Pyd00apr7mgcok/C2LCBTZ9nhER5
9Z4u1YUDx8yAH7NR0lJbheYgFP2YwdANDFnqgh1518CqQJ6uEWPn7TEiF/WCecSP
yBKL2scWN3MThjE9mifukSucmMILgI0PU6gEayQdxWVvmcFANyiPGGLR0D6ylH66
8BhBvDTjG4f9yUYT+82ORIsRtYrcRC7bEfNHsxRk0arlD69NcSygrIXVSm12Louh
iYO4hrEmoUl1Ztv8uakPaVui8EvMx4H8MbtswmS9hv8OQApyyYF5py08i+3tu/J2
qIdZu6Sx0Q/gBTwhm+wYI908TM6wzfsJKwwtJDO4rU2qsH6Ff89hlJYEu/0LR4LD
g8dv5DqvJqpdeq2GqAVNEQsn0BwcfzKkVt3ovuorQwZc67zIFJb+bT3A2E+/3Y3I
YcNpiTg4wuyBHnmeeND1UuooAcHjRkipcb6KdLBq2UErZzySXeU2bYloOrAoy3ip
M66PpLxIXb+0u+FZR7HQSXVYVpaf71Di9XIDeor2p064FEq7jNV9UuBbQPh7cSRy
A4pyRxg2h7/56ck2JHGjkVcS2brrYh14w0ixUCfMUbGt2NpFpvtv2S6r9TJuNn2D
x37mUmmvKMoEbN+HH0GH0BAlcAMiJ9SMEl7bzKGKPF6hylmo0wXuDY7y8cT92bCv
SjnCOj23BOkPW5xKSiAa/2COWhF8dTVOyKtQsbxeYk5evaNOwF7T/mGR62kp8vv0
jXBawYPgMY1weE0m0EZwjXcxZo6m9RceI8PC2FIN8a/ckvlWT9J2vjU8j3h1qkIz
AVPiwoF+LKmdgv4V7RBznmDluX+1kpiM6hJMLfGBJh0phGF+LNUGdKr2800uZQEE
9VYy3A8oNCI8yt7CKGVGCtw6e9jLSD/CEw3xSh9js5YjDLtJbkhHNk50mqnrXqp7
3hB3AxHiWDmmf+JCFCZKBKNp8+lsiMxTJjPN6DxFg0+6om4yF/O9s5rl0bHI04/y
wYMfJOApJsUXPJKOTZsDQxPH2412hDW9bGg9jHNkrxrCKtKyUfSXAPaOAWzkN7ae
cCoV9IJMhZ1QAZiGaOZLzXrsN/CwXjAlrtOrSp5LiljglW/dyWGG5x4F7hyOSLqc
SnufHfLV9oSfd84UJkwO6D+hHs8tcTBhzmBg8JVJ+D4Re8gdHZgm+oLncOWKbj5c
xbFMj/85ZmQtT9hryhtfSIIW/DT+L355B9tQKFHIHncaxfRrKMPFqmIIyY3wc9n4
d4uyE4nBq1CL84XbfMLKC+18UdO5IPn5YFH4UerSrJeRN9m/gXnLjsYBVDWYWCep
wSo9R5co08kjkdOpYhgv/JwPNu4twc36bqaVbKnVuiQWVElmSjZnCGjki5BOnhmM
w/kh8DhbxhMB85ZYgMNBeltBPVr4eHxXoL05ht8YZRM8cHdyoji0nRiHcAJ6oN+k
f9vrclJZ5nQPMRe2813MzRptcKDwQn5E6V5FHfJnK0GjQmfAu5K/S2m3EQ0IoQq2
4cP1N4OxsR9AJOrAom8se222cZqBrr39lONICWdWPGUBZpJqBlgfLMlwkd/VBEUw
H0fMfgOjCp8V8V8A9LtF2IIYP66ZkgZY/W5jJ/iafwIiLfQpVR9esxTZ7DFc42Ke
/NGUNgZdDVjwV+EiivPDye6oRX77hrK8rRrB/fG1CLDRd7tC8ZY7HWY2nuX4WolV
BVZ74CRMnn+1xAd2Yy3b/yud6rXaQSbvlX8q0RQDA8Gylt73NXmnjIQZANvXzJzM
EBGELREb+gHPBtHtZ9GNHtfYquArDRbAAguqyzaQtzvikdN8i95MdfXgvBdhYyx0
ps8oS2IOXc3ihybG6UBFzP0kPt+GRtxqpScVNeYg4PKWG+4VKdGUL+lg4tJxn0DQ
PGuZDVZhDwc0APMCooAkrvRpDVS50kLZc8bGCbxMdIm4r15XcGIbCoLssxUj5Izw
uOQFQ5QMiP0A9vMKwcrYeiJpFPbIIm4wjAwKcj/XLrYA3wFKKun/++QTwWN6llT6
6vWJySlNqk70+z8vBswAjQQ3O9r5UZ6ZUtAzYBi8sI1FGqzCwFLm9xSxA7SNnGX8
U2Gok0qR96Z+hjQmX+sfq4SOcLHS4TB+OWPxaGYYRYV0PrM7MGPoQyIVp3Xeqp+3
Sav8irIjJ99J+XUZAPz+XslkHOQ22c2LnBz93oco7zdh9FGatVQFEiFTCC4p2cOM
hpeERk03WgugkBpdmTpgrpHDMip0/78Tu4RxT7TUZG0g5km2gd8bfshXZaEHdhTu
Ee1/FKOU8Uj1FIXGML427iDga3XJjg/KhVpPbIo2ZYh/oHiU9yK5BmDI+P+A/f/a
KU6omJZkMUisN9pb1noO5J8dK//rZhS9RyxpgnCpxO2FQXau1Esqq2EsTsH7WCds
87Jh8D8nrNU6/Z1P+UggnfVieRaP6gt7iKhR01u7I8WvmwwHYQ+99eIfh6PDtnIm
XrBr9OPQ3NkbPThh/04nnOAqOyqi8DQXuyo+FWlnQ4aEelOjymdKHR31sg0gzLsZ
OlQTB8Gmc8yUYFor+KNxdefXYioElNlaY/98iFs2gv2pwaKAdDgvDNdbFzYMBwIy
PGeW2ci8NJhBO/b/pp7AQ6HBXsCVPAy6hef+QwUOg9Xkzxqa3s2AuEYUrvLGwOKN
Wzz/TrK7N9bkE0vvmuTt75hxAb+U2d6YwgwXPB7fE+e3UIyOLxpocm9fY/H4zlzn
Zg8Fsi3Ivqr38QhnK3sZsrUZTJdMkwkWFEYFiQmzp0Cq63GgOFpRQfO5Bd1brOaP
baK8T+c5dE9iMI3pxQGd7+cXzgEYLPfrhLzE6mC78goctSjLNFAy5rkwtrMG/2VU
2porVn15cbeJTaQnADbdLjdaRBi1M2/9uPdVdjf+Haz9UL0j8BpP/pud9PrQoGG9
CAgxIPgqmXEVKmNhLn/u/h5ZszfkJIs0ChfnFHhBnZRSlc1EHxQ7W2KPlZm+pYaM
ocALIUs3Wri/+5WXh1VFh5YCHaxFd8vQcuBRFmvI0pFI7sKjAH4UTl3Dm+s7fkEo
lNN2VQ6kNGC1qPd+lqAsJq8xvi9rIcUupHKTAIa7bnd0Vnq1WMxIEF2DG4rU9XBq
i4LeNiMaP9FzoHhpx560udOEqpmft20Yx8N4/EyrED5I5DnW4G8SQZK8LC8AsXE9
6j64x+oM8qDoxROy5x3nSSPUjjCuYM7HOFiH0p8sS1XUKCjFolXOzl5VzpMcV0S4
xlq6hKovH1tpABuTjEnFbRWTP87mfwEH28NDGJroH01uGmbrkl9ccTZfoajGEExD
sy6zchYANPNTENm/k/MppUoXGqnpftkTe7bcvNyXTZLv85diMIKHvIgMVLZtilGW
XnoQ8XIraY2MC4/FtPuVGmTtihRksG0Ubzg3yFgO7le2xmYUSmjtFpTb4jaDVsav
x+yeJDT8om0fj7zcvJWsSBx5DluHk0Q3EKK9Rw/3XzmEriXMsB+tzTZohjtQxTPa
JMpi/KpI2U1+bXIM0cixi8YhsOxmIfTuuWl5ocfQYQlKiovMqlxtVb5JmJTqPo6V
CwvLfVTRXIFOYpVYivSnQy3cluj+fn5IxHUud72CQjHhBdGW9WX13m7QYoH2RTGw
pSRZcIKR/+YhDhxZnSxMv3uoL2EelTP6hplc51D49N/FlSIot3YtOXZhJaYaudEw
gChtM1+eNS8ddTrPuzoFT1+YtPME+WL/BCxoSpLZk8MoxP2L9Oa0doMjiLY3d79l
ku2YfE5pu5KTFBez7fqwWb/vNr4rc/REwpoEcF+Pe4OIKuqg4aZb5gvpbWs3IVtU
2RrG7NIRy3qdqoKXwNLykrXynz6CpoB5K1nb+NhI4WG0zahl65L6ncjouBXiwUW9
7UXwwD9WsDaMDzzrX73sORsKFLu27FYcXUpUaO0wHDgeZqf+kwZTccb2ilcyNM7V
hLLNaxEL3pil9MOKHxadoSHo4zbVD5yP3NqT3I3MKjSFtco3EHHQYFWWxTN93Tus
Ao7mN+rw0ORzBhq5Xzjky/Jmctkd+M2PgV9W1McfAYMM4Nfz0ZD15qOZuyzg1T9h
njj4L0UEUBYj0yksQxVlo+2rO3MPL8McdhrXB6ZT5xCfF1buoY4OFL5LuE1Sf9cv
im9dn2aSKj5wfFXhaYsFeA6I3mL9qYlk0ATI+cF7mvKNkegqP1eK5cVSs3M0OLoY
Za6qxi5nhlguRUNC7eJqftb6ZqmOkciXFq1Mn7eGaQ9PLblZd5kMWxp6ju5gRowl
On1XnunIx20BSOO0DY6iJamAtwgIeaPbUSE3rjwXgtRrzQphJHtERx0I6efCP/Rp
9+UFCSFBDl/+SOYmnPyhLDM0W+rErHMPHVR7xHlDuTXVwYKLMmwdzpaoD3EwrmXO
PTLXQQ+bp1+zkdap/93+QsbUrFLDwrpRoK055c/a1xYUv6oyiEPjmW1kIZfExKee
PxTn5qaCzP9eY+oYtGSO3jhUKJJBuJWSIr7Ld9UlWxIvNdBMvDqaRk8xoP26dILZ
vuGZOyO2ryssC/RG8ix29oSwsTwyUD84k6Krl7fkEHW281P/RSvt3oZhltnhDO/C
eym1b3md2n9Mk8nRlCl11JI8n5p85FztTlXeVGLqbKIjxzfNj6n9XwSrB++YwJ8H
NmQPEvmo/YVWCtrSbIenCo7hZrgAG6Cv5+w70munljmcucqOqtlwODnSKre0IR84
wV2S7j9tNEKaPZkiTFqyIIrLIFd6uQalGLbnSeS0KvotRGobOm6KOg1zeUCBGFve
ZZeG4CXsi/Lsu5iI9O3Su+fL6nL2bRFyR9mRxI6GHX//uu24wwHjDRCZQWjziF33
OXGGCuCMR0NRX7vayLQ4drOlL+MiTlS6Mg+AxRcZ6jQpmNrykonRr2fh1Aht3woW
y6kOV1X4LOV8Zso1QAvKUT6IhA56CjK0pWXca7Zo0brc0/V3mg5tdEwcKDvmzHM+
tjTwCxyr9g0axg3V9ZfLs/Ef82gO1tHAj6PYPsuRcZW7fChD+uZbtCy8uwSJnEpM
m7CyKT0fbF1T8fC8L6nOtG66LF3SO1m3AkIqiQ3SPDUleGr+J5cf+8Ec+xsTJ0A8
ydhRQfNra7dzMvkokbAtYttWUuNzjwqkKDmXLMN53rvVBKm4RjnpW8jDWIqhrDef
9BiB0rlaNknRmgX+LlGU6u2wvu6eIILj7fvsVxBuNKhnQ1q6tnY7CJhRzbgKKQpy
mp1V4/xZGQXvXlFauugRph31bbNqiV5lERDXaKUfGvrDAB+WN6bs+p6cg1JaLGM7
wia3yOBJp1XsHPzzJAp+sFBpeMeaYiE80oJ0ZALguSVro2SFDzlze+f/IRMtn9A5
M1kWq6KwkJbC+2mCqu+74wBLDh66BjoHB/yXO181euZcoEvTc+8PcJEej15ODRcy
Grt2IkCpDJcYI/t3aVRtI4wlyBgxPoy/HdXUIakv/kFwVnTgwCH5MECjzktRd9+0
SgLMIOfxjHAt71gSRno2xTxhPq8z/gWO/cevCOOD1mmMsUIeFsd9vM0Z6pDaxJEv
ZNDQ8p3I1M2ott+N7Qq8FUCURP+E0adsxTCdDtR0/uf+P91tRaiaZNxYthN8FtbG
IpK5ykrjfxCDSsV1d/Ge/muzr03yHShCfXdadFhzeJvIjTuQX6NW1QrxsxB3tVca
iZsc69K7dwn9gAz9WmarnCp2Pix0HFeJ5Y7DBn3UbHem5VWd0Q+9orVQbRDU/wG9
f8SwC+62r7YV5LaEKW779Nn9yvElY2YIlqam8z5fYNTQSiaJtdFTfpwG+RWAAFdP
ViYM9Ke97vFXtWKt5yy1XfoMdwBbl1jtrq+ESqGJhOqUPmtPCDA2+RxDBPeyOH6X
Wjm2LSwwnYMpyfw2V/OpAfDhDds+sXaseO5QbunvotBVJ3VVhNhMbK4c7hkeVQxa
9apfZSOBVlA6yvgmE2WTNYAvZj+X3ojkKyZeTMKi7GznGD88+k70dpBApsvDAtzq
o2nGgp7yrdw+bWQhlJ9fkc+TIegMp4c0IXA2C0De2ToPaw97MaSR3whg71vMQ3pi
VCwdiEhASImuHEpfORG0Xc4vljL4u40CoKbEh6i2U/t9LSoHvZY/zIVMAh0T5wIv
o+Fa1zadiMU4OdLXraEL5p32KqWuIES79U/ptFNAoAxIqCy2mtXURE7b3yW1s8tG
mkrvXyH0gybNFYImPB9CptQmyxIHAcNiXL/a7rZ2cRv4BekHkbo/nbsjKhaSgKSF
pDXaEuLIpyFIWkqWQ9NgAtGoBFEfL9B1+cDgvBmUV5sjm6lPPVknonRJjr+tB44k
z+cgyIxol8GQCGC3RKINmFJzVUY/hUWzgz3cp5OWUfcELKE+UB70daEU+QRMid8k
TACDgxY+SXyLVyBlD3QmXqlCKe93MvBNOADDSb/wcTK3sUztdhkr5bev6VMbzLij
AntfbKQwQfoyciZ980ja0RMJnFUlR+LoUis2WaQBWXvBmmUpMHjQMHaj9RIiu4yp
CTgqmfDiTGlo3BQJu2GkO2pT6nZAjnWD4fCkQg7k8srlp1w+GvWSfBPPuYGLXjs2
RJzP2xYk0Yvs3ghgqNPZoQDjckPrNR3hiEY6TKkU1c3dlePfu0WokYclxYg66Z+r
MbNtUGfSQpJ2yCUP7U7e8DrHa2orKI+ukc3k7pehPqTBxCgFBhGiCmkOVkjntdLR
xITDiCUYjkWcEqN2TlyWmkegiJgqBejnbmFlhgy2By+JBj3IhDlTYl/DqRAjRD1A
fmlbzp7qX0l1+Ei6wtF9HM6HE87EfQuhymuVCwFN3t0Oo8GUZXUXEi9aOUwOp4JJ
2woQUXATJEvRP9mUR7D+Jy19fjiA7UvWDtKiYCb879i0e7ooS4utVGn/BX3xK9v1
Kv1/1wRl+xPaJ3lcmwxeUhagyhxQ86gKOUtyV157iLXKTP5hXnusRuJatzlpEKpx
n033hmlnB0vJHoZG8dziD1++jmhU5qwDzIqjxVXIzS6Z34lb9ThhgvpgXTl5p2WK
Apcp4DQZItGLeEVnAH6b/utr59vcfLv9Q/OIwqq//NhalkCd7c5Wrso9r22JoYsi
La7OytfHRzYQbX2IdmKfukJC1RPneeAE2DQtARwGcJIhiQWvFMkvlInCNb4/nL6H
8/LtuztwKmifdHbacZUWHu03yt0+G5NvlwoUEm7uB4lywWszJSLqEZgDQMdssN1G
2EkjaYDezJlgTgi52JgsZy66P57sWqMYfIxxTWC7RHl0JBUpS5uP7Q0/l1RG35zK
LvBe9XrKaPCs6SzthujHZf/rde0UztGCgiCrtvtESK45PlYksaLcv///2oxxDRVn
TsZ2EyHLHN3ap1QI+UmnVZrdeq6t6uAwSdc+DK+ge339pJ2EFdd5ytg8ZHy1oKzK
2Wmsot7ZSqPOZC0m1x6qPpsZTRBRhEoh/bOTHdwpxckXGcevSCAHWMMAf85t9ZI1
A2WtwensJonGQDGI0LiA0hveqEOI5BVTB3eGqIrQKmhoZb9R9sKHCNbQD1SBEi7H
xgxyOv7Klzr7qlhdFiToLJE6GkU53aDD1Oc3gZI+htGyG6E/Vvy6qglzL83oDbFN
tsrJlL6KWCtLofVQixWw6c2z5ajsA2BU2FSXTpGPJTk7IJJ1Q4dSj/+VV1BxvVXl
nDU9tsYed8AvX90f8W6DM5XkA+eJ1J+YA32h2Y3e4N8kfCERxByRGEZUlEKnQgDx
umJXJAoyKGHd4p0bdiyzD4WxOYMrpdlkVDo85rVC6PtH/Y/A4z/usmheD6R9OaOc
bLVeVWqyXBnluJnhCCRUHYzvWkq/Xv5wX2C3G/+jq248HKTgKEKBHo8mlkb4WeL9
WYWzhKYpoHE1Dg55+zWJVxCFXRLBl+6H8BgGwZ6MIw655HJHHJ+4/KwiPzew2EH+
H9IkoP8qU4rzJf0h6KUhHp8QUFNcfOgYPrkuRSbE6yKR0J3CLWmBFTwQe/ADPS+6
5QDg4FxC+iBLLv/C3CtNmVPrWfxi2lMFYjS+HRFlqXjSuH4k3ONZrmky3o0CeeG3
xzVVzWKf898h/SFrzmsthF3AGnXW+5zpor/IbMzqX6Do8zvRA/qUbjB0mElWArn6
wTS/jzexdiWh0ayldTfYDeg5YCeBrlKKX+ATBkgtrjJd0KZqX8CrlRO/8OUXkbd/
PPoLe2tmtSVc+TV3Oo84KbQ3Wljwif6W+X6v8JzVyGwhxMCfeF0obo02B2WkOZ26
tJNb7muO5MkuXIYFkwvitxsav5ad9o9xjYFWqleDFzxbHG30CFeHMTJWDjYLA/jh
JIyUT48cOQXJuZ/7kGVxAB5C/VgdnGEnnugFsoeXr8rqQCfh4lWYDNkvw/nR0cyJ
sqQ9hEF2/G2AaAAu2PtbC5mEbWWB112g5lLdGu2O/uXe1386Zer+nbbD6ScIKU8Q
0uty+xMibmLDPENzbuQU+0LbOqtvFVoYaP0B0afk6Z9G/PuBDjzko2bplTIgtfO1
94LukRRbIAI8P5oJzLSKcCvSAGMMncfZ/Vz3W3IypHb/4RNcnVT7+UdApIibIbKI
rgAp84jRhMelnMHJ4iK5V4wWtLnHIWz2U4vERYDic/rwxOUYEQLZqOdzN1swy+0D
hZvk7jEnfpwnlcl2OrZ+uDrywJTIWfWDAzYGCOq3Bin33UkRJGA0Z6yoS37cYVmt
rm7280ghRDqdkCZn3X7K+xVjFrbrvLytwT/orG5I9rYsvqJSzaWfCg36Fa6OPAK+
/xS44baN/G4PdL0qbw9qsbDlxQGVNC0+CHXL/nj2VkZlySek+fgLDTVAYCH98bj+
YN87tsQK1hrCyh3MdwwY81F4J9bJZYdJj3mKEg2IO6Zx1jbPGmD34DbGGB9Xbq0I
EIbPXEXG1xmRWoN0oPGkBZi7HcJ3ag2MXUfkHWP2FEX0/ere2hksPk/xPRQqFmi7
eV53n4LQdKM3rWnsDCvFCZs6O8Z4rHIVlEIqhIfCGVpWRP9XJFJcdtEm5e5QTgT5
BDqXNE39k+sFvVKqY6i5RuEKjyzqjBw0prD9jsoZH7XlluzLD/6J2zMCwQ9VHqZ6
d/zJrP16xmuO+zoe6WvNKHTe4ABl/eQuhHC4kJ7wvf1Tl6WaNc29tddEwOw9qiLS
MRlJAwlqihoykkMqJrdXB7yihVHhRyOy9MZsFLsOdkDfvjdqIqe6yRUqJSolCznK
2gTxdxsjGBHhRg8rm0sSg9C1h6tyWDoOmKA18lUeL9AfISSOqTUcazussWqt6qyI
jMvZ+RuFRh27kWx1IoM/7MTmTarEc+xzt1gJX2tlOv0aNyGMSCfPf0wIBFRTcTe3
hwI9ttxOfpWG9iDNaQZj+PpUOYDX86Msdm4JK2R0aixFP30vp4NsLp67NxZSOuhc
Z6qEDYXZ4jyK2Sg3t8NwwGn9I6QKdKLRuQXwVDVYH3LqwZqoz5n39xXkeimeNIlt
VMDc9w7Ej5p/bgokxsvD8mN3jZAlcghvr0kYaMasj9mESE4hTJS0dImNeKbCw8kp
prkGSU/2OrvyZMa9bMmtzYgUoiGUoM4fQ7PBG3CIJf4Yw7oswp7+dwZLwlL1bfkS
zVGXJAUNaQ2RIhucOhwR+BcN6kuQy0acX1Z+MMF9IU8ouSmEnlr/+eST0/Jveo1m
hZF4/kpOJ9eThbKgWKVGpNulfdRzEMjkmaAQlx7Qe5FdcjPekowgQY/tKMtQh+v8
F+Yg47hjk98ljK+Q+uSz+TMz1iwxJ4Wdfd2CJRxDCgl88YDCCa1jvsW1mUrHwcqH
NoyaH9+VUcWTs/L5yxvkZT6uFqS3e0twI1FScHIMUUdQOnvYdcns50WoVGq+JLWP
xJc2JtODnZ9xeEFsV7W4L0C1NABS85bAFhX7W83P5cvhZJUTpxriGAk3JDMpXIi5
MJlzP5DWv8qzKGdxpK7eNMX7eyMfGTOfHqUd2Ke5S/F9pyvIcMXoo/Ws+MfiF32C
sR/AKR9bGA6xHZyCpQdjwOFAUfTFbviKlH9OxrOoxgWSdi99N4eE5PVobwRxVFrm
MQFC8DGFe1Go8dYk1SuH5kpMuwPgJ4C9DuMgnCjV9OzLdg6ETxUZ4I53bDDIrqnh
50kV/v2d0Ix6G0142jBq8Qr4RaPiXrzT9ZnD/1dkLy9rA20P5wAHPSnbI0KdbKV+
ZfSMm+V6r7k0/9ydnFES3gUvHDJBh2Cf7FnbXq5y1+br7Q/EzrqvFZy8pI+IWcIK
Kr1BznYf4yHlfxAq04PcLABivsi3gg5nXcs/Hh8tck76oEfnJ+33xnCWAl2TgS2g
Vetndsir96lYNLAliSpTsdZATbw3j4oDyrcqGenTlbyG3WiE9sSIMKFoK3EkZFy1
Lo2F1OdCN773JldH6rv7FSI0VYyQj4z/xv0Rm446SIX5F5tnm5lOIDR9r2uJM3f6
OGMnlVvltikZo/jtoUeufHTxpwnH0b+l54rNrcxcXwWU/RT9RhCkH64UDP60pDz5
qcNOvEscNcQ/eOQj+r3zaNGUvWPB2WkpL0TKDxPNw9cG4irYU+h7hW4ETjMqt0VS
W17hKc/wUwwiebf3qHH9p4yhZvWdZPz3avZPBoZP5XG2togLn1aNbB7+GntsIuY3
CUqIH4VVVm4tKj/sX6R+iHEaATGkPl64Eg2s6r7NkceFvB0+7yq4pVhRf92YQeZM
XfnOsUwapp3IbOWkojyCKpvbl6Ts3G68hawrd7mGXXNs9ThUaJrVwXlJmSyICweZ
0dTUIkN7LhrIQAxocdPYpSU/BiaVOzZbaYvaD9LtfjjgAu6rBuJZsGw2hWWWLEi5
2LHfRyjgmvURlGQT23toWmw/ZsUnKkL6u7Ie1WD9VAuWqqJ50uJIMogRbQuQ8lyh
q8zuL5uNuNYs75Dh2y1gQBU61qwtPYt0cGSTgAnxQG4gPQOVrg/g0T5gtHR39xfJ
386RIOI/mj++9B6Ja6e23q8B1CVy/Kpm6Zv2a9ZlMGo6AyMcJyohBm9Rdlng0kgt
0fgTaj/Dt6AgigHWMVWXBo604qwq6eY+GB7UJ8QnRAvHsZqoT3sSOKkgdmGo9h4R
2qXQX/E4vPRjTCew3xxlgP76O7XbCrS8snxHMvQRV2qZxlSZRHXPtp2eTzHDf8Ez
0e1n5D7dhu4Qi2kex2Gj/4KtGQIuVXCSo24BxYtM4vwdvFi6Z+5yO2dFYMKWikA8
bs7KTgil3eEOj0aScpn9CkE/skruQ5MeQ9Vfq6nxszxoCByKFhzuKeBsIsVyEdY5
S1Vi/rc/rVPYKgy03qIaijX1eXOaChTABNiN/eiL+h4WH3CSHgOHG8Wdopj7cc/z
XE+CrfcmAoR4CxCH5SyuoKfAkcTjQvtFJVHCIduZ5VHKgaIQV5/yUD8RVTFtgMl9
4DyUuPCsbQ9An4OV0HRRp808BN4smhugP1PAe7Mtwl2Qz9yd83JgOIAiR7uqoA+g
CX2hKdy0B2pwxUCCXcjsQYQaYjnNfBga+fFyPY/6RleJmARWa5EvbHjkUDxTAkNh
2AF5m+RzWnfbSo74TwYE7rndDi1kQ3+vD3TjS+m22NPqriAHZCSUVzyt2AdQK20A
3l3eEoY7wpMi6zS3cUeRE+IxWnUxCrfivjEIF0xmVRgr38pAVGBquMJuZkraRJKe
YsfuzH85JATTrFShGCIqeTLNvu7wu29c8iBIu9B35pQvXqHkrvnYPseQBiVJw47m
gZm1dV+OoZ23DNFDqsO/fZB5nKtjrzm1u8EwcJfRQYu9J449y4QyYWv4fNrg9kUr
1l8Eos7OYssCbz7Pqf5ox3ye0+OxKMjKW4eFVxFe2H2wGZBu+x9MudAykDePPKOF
X/H/bE2D2wsS5vbe0wkQb5te7NgXSBgYqWnGFBXNJcQqw39mAlfz2o/rdf8uzvjA
10k0jyo1o8gH0WsDUUgbx3yqiF8+E2PU2CgYEM9Pi83bVcHCkoHqLxwG8z43Ttwy
+lX71yX1tDIMlYBuk0roAR/ULr4SUuGDikn7kPeQGavDD7r/50VdXFzm/JgYCTZx
y4+Bvc1a2jInOxZ+j5sXWdumlXST27IFeyGnAlzeUYMlQplGZ0gb1lc/54YUOEJO
Z1y2cqd7msuheCwE7VCzk99csG6ChddpO/XBf/TNHsze+jUhF3f3vJRvxeNK2HJ1
92LK8hCbkop2CM8EuYn5tYs5/RJ49eHIB3MxWGkEcYLCvorTXF8O9EWUHTd3nfHe
iQ9Z3FT6Ro35pGhRmOKDUyUea2lVKWrnEtsUQWHN00tmcqFn1QSSAf8chAhLi1zH
6pMP1c9AiTFbMmb+yzKAD94M1TSOxne/6Fcc7vicsOvxm9warslGzagAUdhhkSrY
t0TXSMKXzPXzo9pXDXEXrwyfGa1E5siN8bPJVFVxuDNtjTDa/R8ex9UjwEkiI/T5
dE4JWo9hT9YQ4HbJkoepkUdN3PA40hImPN3JOtdSpLJWq1ktHTovdgmrDjU8OmX0
P3Bd7+7kAN6oJRHPJvBq6HDleTSNF+aZZJ4TDQ+yQTS30krNhmfsoaAMY1+CSufx
JfTaqokahoBCE70DPWt0IFfr0Y28x6ias/aKRsTURfOfDdhgM91+7ygpmfbqxNDi
focZQ/AVP4PgSaawl6hPj9w13z5EMkhCwyK4SeKroyh6eiT0pXLqBX38tKvPQ7aa
YKLbSTDdRYCgHu8BuROTEuOlI1MJmax8nmjrnuB3XM2VzSdakwnATabuOnWI51ml
Bqh0YbYJSKd/d2aNOEdXB2/52Vx678fm07D3XRtIJg27LUo2TnmgLPgfALGFZsdb
RYj4Ql+EXmvdfLH5fnpUUqiWETonxmr7piIMDOAY7LaYDVkztB1Q6foSNmP9lmTP
aMtpbdySbf6GetX9UZICnpRLtw3ge+Wuk7Rf+JHdkoxGIXH/2LWLn1tPMmclDaoW
L6iY/IhUki5rVK9MkcXAVt1KGXZZLmSAbvljKwkKanC3IbdUxsB+CalTc5zrVcCi
NPmo/jZa8E6mwDo4kOYS8IQFbKu+4SzQySY/x3HgkpZcpRhi3KMfEO7Ddfok2NFk
X5yFQDUugXeDxzXMacIALD2C77qMraVlbKjXHW6aqGxhmNKW//VM0ALhHn04qdOF
vupCxKBZVhZQi/Wd9RvBn9qTFG9AkmXp5D2bQ1VzMRZWq/61wUxgtrHeBX78CFCy
RcpRnDB3qMtLvTGkaaKUYCL4SNYJyodQwrHbrPA/wiK03Gb4B/MoNuYjfhM6bcRx
u9+p90TdA5+O+hxFTHWrNSj83nCoO9Ycq+GVoqkfvSVil93cefw8CDBwfDsdd8Qq
yHbCM20inunB5QUSwymFhX5VD7itpb1Xicy9qpOu6OGdA/xpuAIIA9s5WjCKqy2Q
ocehU0xeNxXZ/in7ihVUJluUW7RTp3JTufO8/YpTiCjqmGoNb/E7R5btqbCpgaxM
EWaTFoNfc5B7G0AWv0ngH8uz9w3pzq6xJN2/sn1E5mnw3AVahG47231pFfGl2nWU
K7ioMEkGrwIGW9+cz+ytDAjXksn/LSDuBIAy5m4qS78g5T832MkvbXI7aByct6Rx
WzzakLEKrmbJsvP+lzrzWFQxi44Jow4haz+Vm1MptacUvh9oCT2UxH2rZqUDKuFW
VwMCdd0lYZ6UcuHJ7gKHdTsKpLxnvSqR3vXv2xpiSAa9Ln0HYkt15eOKc1Rbde9m
JzQw/k9+E7of0lUgH4DHnrHmHjzTSalqfGdAGTpRpkZDLUCydOac02vOFuVZpwNi
70Fu9hrwge1LCg4xvcRj/SsJa9EhGeD4LHUYavhumIE64SMASce7enrbmef+whlJ
4nNng3UyWBhZ8ZPkwSRGnOUFTvzqiAYJpP+3MhfGMEStSLyshS3mg+JOJfdh2yE5
883fO2YXB7jTADNa0UAkzhVyEng1WyNtgdrzzB5xWLvW0tTL6CgaaWP0To73r+xh
xJ6EaqgqCZrQfiKvdEohh0UxX4ftGuvGcK45E/9q6CeIDyt2RDsLGqGCDp1KMU+y
vJBL02nh0ztU89e08GdpP+GcRXNXDBv1DkwtAiAyTvNjLhyYzlUgOV3GjVVu1yV1
yyHF/xqhPqE/Rx2g+w3fnO0btJm8C1v9uL9S5nYz/7nNM+AwjhGFEOWn09tBd42g
L8d2m+D6ZMKxZUhSQdnbfkidH3C9QDDK/2R6VJ3SXLSSVu03T5Wxzl3WygGo5RpD
XWfCifIBD922x2zKp6dfT4YxRxhokbhMfzwl/SeTKyK7vggqnUk4PQbs5bfPAJVa
NmgMfNJ0ABnDv/Ay3xm6ck4y/br8EsCWgdW5fLU7yMSGgoW93SGbH0zygsHx4/4C
JPSB5Aj6L+LTXqRTusPXPLjgqOazEMA53KWy/dYKc4rbvGUpjYUkLomqw2Xq4tXC
THshyunNZe/W9OiDxDVC/t/aReEgvz7berks0dqF3RP58pLCskCm8ThoIjdtqKB8
/QXZB0aVEQNmKB0qSDVBLRpC3p/pni6sI9NoABEyQ7+25X2WFQgcK67Jf8UmOr5Z
gywhUDt+ZFTS4JyrARcSHteX0yvbtXHunFycOOt+oHn+uUPtSoVoRmxzatoycuUk
wlBCdt/kE11xws8lKix9LNRU65XAH331xeLrbMhwt2cNHm/UnHyXN4HMeqA+y6qJ
oehmlSCtBugAGEYjnZnAJW8FJqpkaDNNJmJgN5c0KfXcnLNIl848eaOAOhN4SI5Y
k+TcNxjNOegoeDXL8/zF78v0btve40URvTBqkPh7EWMPtj5t7eX6sV0ciL+RddR8
j2G5Bq7cwuA/68/zf3jfWGyiXwJwo/LHNLxqgG4tctsY2NEdCO/yGALfTzpg+4Mw
3uGwcvrrykRYCeYqNrMx5EDUmvx7Y6AnLpW0eExfX45AGxVvm6n34PU7IYI0HnCS
l+5QLzM+Oiyd9dCJGdcBuKyU6uO1S0hhuzU85lsIGjtq7KzfForc9ZlBta3Tc/lL
qDeyW/lcGA0U6ud7vEXK3pXzdUf10mp4RSufcnnO4AAA+VASz9ushwjBDlHXQIuo
4Rgdq43GnTvbA2UHyHHBL1f2koedLJaS0e9gvRQq3ux+KnKCCe4P0UH2YjsDuxKV
rbUY46FajPwR7co6VZjBAIQYAw9RTn2L31VFFpjLwexuPZLN4HWy3QBddIounWKv
vbRFjdVjshgj2bSX9urT/nQ9hPF0dKRrHjDk2XhdH1UeooHNsvT0AFIG00PI+FHd
7QH7Uj0wvQuGbJf5ZiA4kn9JhDcr1I0shJi7RuuLAgOrPoEIcpUJgdjmbA8leRH9
YyzrWUrw5II+Tm+QzXDNKBWDSZaTmlEqXfxaYjK0NPZao9PJmQJg4oskrjHS7iFy
HMTkALaKYhsWxSt417C01zhcmBp545XRnSjljHp8Nth9PPnb9dx41HLTwRKpalCm
GnrqyVrAUyFbXo/yKg3toxFGfjNG0bS2e8Js6FFWC7bSEh3QKnL4+USm96UvNRzI
vvhfZ6gDEaDTJdNFva5myW268hTKerVcnWteBWivCVmEMvPAsNetvaBHVryl4e1E
ENTDK7knvVFuX6H9s2LWiAcWdcuemAswpsKQyXV/NdQvL8XBH8NuMjQP6HNQW7id
NWsHLpUN9sQ32GHBpOIsehDNQg3lEjYJo9UKtakiOwdHCJ0atPuITZpj2U6IGQLw
crq1XObki32Z5Frxr2GWK/RGotryH3OiQcPKBjknv/loOg1Fmns1rsanUsP79C0u
v2xBwHs2fXerrGhbqF9VuxKUs/BHwPwtrErQx1+y4+uY25R6wF0+sXMi3Tu2na8D
tfBG/wG9UpGtQ76AMSKXq9+Z9kNvavBBZZdpfziElP/xmCkqWnlOoGBfjTo40Awh
45VxcRdpfY3M7VOhbdoFHoh9gdBiD3ZX9SPiiBpCdaOJt0/wqOWHGzVYS4AvgVKR
NWZmwoBz0ssqLBzFHbDazKMqtO9BHlZHDXM/WjguLT6/AUb77smteAYySfQgpYYa
mn26ygIVtZglU3dhm+5YrgnbchQPAxByyf6FI2ZIL/Cz1G8QLhP+u540pXqPRMvl
bg6DpRPIeXL6+RgjEwYm5aFrv5oMZ5tUajpBskAoSO1RBIQBOTczqrAaDs7JQTJO
/0OqeWIosLNyL3sqtear0l2VB7NxqnYxFr3Ia7+EpQm9B+s03KBJNdf7ws+9cDpZ
rzmHb7f7q1KtfY5WAO3E1u+MbC/d4oBBV84g3UdXHcoJJFqYZC3cod/BcoDcHmfv
HkBhfAxMVyFZk0N4eyYactxgZO2Kn2mZK55ukCwGIA0lDh8Ct1UoGuTFpD0H4TAm
9cJpDdX2PIsb4EveuwpkAuujp9NuLuczv+JkE5sbycWQCUy/ulTumEPjymfKVRf/
RHB2qJlS6adK8TAIHFIQXbaL7kCTYPp5wo+ViAb61EeCCByno0UG22rQp3j2t5P4
y5n059PTqFaafqgsN85BUIBQZWWXPkma1dKQlM5hno0uWpFgXFTpNUH6EabpLneU
GZC61qz5RCN38g6qqs2TwxyULAvKhr1gE4liOiOlkQhTfithHWXQMVcLVcKR2IWG
XFvWsYniRB2njAIEipNXPqvStj2UdVu4VSdqHqHth9qqn1ULmYSWKHJxBut8BzwJ
xakuXOOeS6lMvKeXylE/eXx1VBqi1bvtbwl8A7CthbxRyCTH/FprRQI1tp+cSrZK
MB91jFqPLwkcOCkwjIxaoh9WPmFjPOB5lKY1wEgi4kd59W75X2glJ/kGMJJ2ZZ3v
qNHEae8l/SlaaNWHng2qsekjHg135cJvHH3f8cFBfbcy4Gi0MsOBp7eGfPEo1dXT
3CypPx83fN51a49avti0wV7ksMzczE/o+3BrrjUuayjzFSw5yjMBwhL1nQ9juhPI
f/+RSUi5W5tl32bkWQl+2ZPGQBMHwzjQVRxCBdCMoKABd444YPYcit26L/PyO+mD
ZdPOUD818zfqIpRSlmfAGpn/d7Urv8hRu75tKh/a8QP3OcUepURc/zuaXGDBOahu
4biAvs2lERmp/1FnYAJPhOwtkz44v8ao+h4U5gufGob0SGHsapvkNy0lGx82p+5D
7nqwUsV9bbRLQXoqjnOYZuXCTCH16QNmxAEo9/oB/hRd9L58HZRx7mZhp3MJH6JB
4EjspR+Ka8XdK/V3O/w6OdwprvAFzlzYL5MN8Q+XHKeIzwx4WYSa8JBMfucUFeeD
xnsg1E25xDVfSVy2mF8p2x5+DPe/sGxE/PnuKQUhy4HceR8eL3Ipd8FVfSnCobmc
W4nlCumicHwnXEbK0+e2I+MxxIJyfzUVQqPmNXt8EE+27EjK+eZ3t/xkt9pHno4n
KK2H06uSuOjlYLipiizCkLFpTwfDCfVqbFa9pP/hC6Bxc8zlF+o8uIeesr8xM34M
UMsVohEYKar8tONBgYFED34PHMwCutUrVJ+jg50BQYY6q5supsff6/+uxYp/Xus9
dbTxoxKlUTquU93yyPMzqKS7WdMAgZzT1Jr/XE+XbevjvI2Q9KawrOH2G8vg6PKe
Z+pPUbxzGJCf73x/lfsOedIOqj/TFo1hKuYdICWi4Fi8D+tFW8JBETKYueRbBn9O
3olFhYYDxy3wdr6z4LFaGBm8JxEQxG9v8PH5cLNWNIW82Lrv3YH0gyt5OYGlpHbE
wibRIqlyJSkoKKTeFVCOdw3uMcBWRnMZZSrDpSRzU+uB9pvCQ9ArLKCPz7L0F9Az
Veplhnw8kLBgo3H1PzknVhX5URTIx8BoS0NUKkfhqqggDyu+wYlQiZ8wZTnfVi/3
IQHDmifoGfo3HptLwXZAgKS5xcjWtKJmJKQV0PyhVRv8MTz9E3WgcpyYaPAUOMd7
nY50BxZHfsomlqxbo/y260lmu+b4pUJM/FOQYx0wcY4X3mtk9FAAIk6TlNkg6pO6
HnX6I795PGkbs8qFWTmkD1OhIFJEaj5pyAhACA6k3LvsPEhvN/xo0ygcwJyPgLcu
Q1gGFCntxwcyDkncn09Sg5YfNIhoJmlRXDRIPRsaV1AUQwyX69ouHz+6RGQP/hGk
qMAVh02tBk2uPTXAT5SlfqHtIzqtX9lf2I0httB7FAAoEGNGMzTsah6pVoTDhkIG
qODd39hpdef7OfD96rw/ptsQQuTGYtEsV3nfE1bwUOn4AJmP7K57cNgW5glbek2F
6ie7r6Iu1EadFgCWE+1XuN6RffrBmx2VPH1zHGHnp94jWqFqaIwez57YRhpa+ZBG
6urD9iHX28E9XTWDQQ4+VOD4tn44zyt5FW6BeOA9YMabLiHYQB+yVB2hwFuHWAt+
IL7Hg7nPgxp1bQ9M1VbCFBw5hA4vT7h8w2eAuWjAH4WUz/hniRAm7hDcsSirZpe0
h/ocaAKgRpbPy0VkJiOvW9CjaT69DOyp/5a8s5NA/smwY6K0cHUE2eTlwzuT1oTH
dUvsOTBfPk6tzZyQ502ZwfIJTiq2EaSAFK9xpRCJEt1t7/IiuvOVBwnReAWNXwm7
Q3vHo/pvzUW6uiczFhK2PaE2AtiqqI40ioB8PSvLtYvbdD7nSgqyUwW5FStkKxuv
ADIWKi7y1RutGWtncw3gz3w5wdFzVVWJK9C+q0fBweJeWDtM62iZGu3vTSkVNuaU
UZDHO2fowSPE2ldJt2t+uiVQNCoIrn8HHH7czcUde81V4Ysol1u/iSKuLBBX9apq
uFrntMK8xLvczl76lrtGCYmuRbQgAwhBNvqOvPCvRs3qakgpj7197RP9VCtaCqqy
sOssQNOmKDsxsvVKRqdJlGCKXNtk0+5V1dLdxTz6srXnHK3p8++pLvBeOodkTQlM
TtQqT0283gJfsonzEb3k2IOACUl75380ZQjqMsmzdOoQP5FFu2dRk/vtWwLb+APk
qh+CYr86yjOuZpX6+kNHgZyFi6gClejiFDN7TN2C6tn8KtIyLtMBMS6BMMsO8Gfs
kgCgoI60fQq0qkjSW9qyP5EySjlooJMcm1L+bXFufDxNre89PJVA5AUnRf+qHLG1
1kk0tnIqRbnob3nZVjbdiY7SatpJEKvzary1cDR0PJw/go2ZOGZlIoUShtL+TQXX
GYrDHtErVkmhl2wCV90l6jirFdoA7oSZ9Glg0r381pw4Y0YvueFTkK8LMSBJ6oX+
6YYZ4lXFy4PjxKgQry0DkKCdmaJD6CUS386h29qoDyElI4ESjo4VTTmoeTzN1qYr
iMzPKUgoMAxQnS6qsT4wkfBfsQX7TbTdnCND4eW1yN+KLTHKMK9oIk8OcmD1ktod
sC3rmyuGRM8WUASJQoTq3cFj9vdgVMl9P1fZE2Bwa3EuXTUuRmOYvP0cmkWzlS2s
3YEGbOdZ3XBhELlMJKwhuT34xeVzmhbJZMnh2f9SEkjlko6sWnuBPJ9kmd07mXnK
Z16SnHUhZgO7/rH8aTRYpO4zqEZyuly9l0LLZ6q/iugLqfhPLCWDqazPhReFE+Yg
g2wMMUAjwP8BoeW3WiNf5fTC1cr/kVlw+IisxG8ipfIZ6mSbm5Tb+/191kx/3MtA
L2ygO/GzxDtxWcnwz6pOai2oEsGSa3ODsGQuc+l00jjzsfSLDRMSAzWUudiczBC3
8JscvmgZCbfzJE2+ji+23RNOOm8uf2AUZusuryPwxizJe4K4AsAQGdJhVOOXqqAj
ckFjTY5sHL/pKkFapAnIVZdkty2ZMFIooIftsg3S4VmJDVBImXYeu/JVR/NxD0M8
CvfBFOQ7RaC4SVqGUPmZjjlFkyGcTpcvREms70ivsxBVJ22TfBLCN2IMaB4Pm4m5
oWTSTiUkGg5P1RFFzq/1WQ5/dKh1A1/JVBtn+xXYVyWb9bCP2nOjc+4MPHOoDHOD
fZXnEZUhgdacdmxS0TWvmEtqU7ofz3zn0H5NYiAGRPLx2H56LBtxyQMjTjTrXfSP
Ba4qsR1naD7IHKziKOFBqvLtiYeZgLHdMyC8wuF6T1ZKSx7jY/5KzhB+zzCscfJM
BmvIGIs6eFrbZHOW1PQnR+b+ovIGVZZBNJI2gnLo9Ulq5mcohMZvyVga9XTW8Akc
7q1M1ttMQ3lRacVEVylD5eNrxj9v/II+9r/ckj6Bk6h5wvyXh8eUzApbsyuldfcu
lcq+A8OPy5HFPWaCF6JbIJOt3b6nNpb/hy1pClBRJEqzzujytCzz0a/nkqN77lZE
s6ClsaDe/etzKuhpZm0P39xDY+G3L3kyp6xckOH/88S6fWOTDrrYMtjksJ/7GMEv
fWTW4wVtlILa1xxCDphKw2CW2iIZtRq4XW1avwdilT6QtUs10w1tqGbnhxrvKHWD
vfSeGnqxMeztTPAKEbUyzpCRIKQbpEO3p4GooPijC1LxHPr+u6xNPM8H1yVcfZ+s
thUhsqyaykgMa0bPatWUVV03MkBz0b8ifSQK7uNPUZInu6gxx/yHdrEC4GZAYtKg
V+g+mAZuwU1FbXgjXueoiglpt87zTRC5NMoFgSsmAC1Swjt3bNg5bPHO4iwqzzpy
ZP2w67lPv8zKu3tyL5KcO72/uWkNq6ro/g9LEa6ErcdsLyjZz/zuS07bKvi/fvYp
dbUpxG0wF9Ocu1PUmYCxNC+DY7eU9YEs7/zUPVo8TfO/zbkE67Cf+VOf155GKBEq
XPPhJ/IU9t9eVdbwGcX7ZDoV25ktKbuGaEr+xYqbpK/oFBA4AvroWuC1U3lOuUmH
`pragma protect end_protected
