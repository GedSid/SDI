// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:43 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jKbhvdQTFxIbyAvRbilhjwZ5LcYt/nErD4uF/hxVWHdDCUyVnR7B/koERfhapQBQ
SweJcqO+1mpdz/EZEWi2xrFN9kWq2ooEDSXacx1p1wTsKXVgPp11EE0EMkaP4PBM
8iDs5qdUVACTwweQDHw2QDzTSwAcW/U6v8jNHNa4r1c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2288)
SbmTq19XImiiSDgGuw/tjBXxNvmSd+Z1mLaOuYgyJ2JGXmJbH/PyNoyd4zj6UER3
/XH9VXYkr/71B3Y9A2qtlgzT1/g1bp9uG26seyQ1M59xb3MvnNwS00/PblUXdiKB
RJhzPlnibMqWkXUKF7xeY/Ub3+rbIW8xtNbIcFpaY4z4f+sA/kW3OTokkqo1yDWW
vQuE/XQ+F0Jcw36+ZKiIeYurmkJbwBbAcVzM1PuKmaIAfPB+Gjci/Esj5jhELTmn
6Now79QcrAftDv1+S3A8THA5RnZiPSZdizRa83zUgxp4NMwPlXEiGzALRIfT0KRW
VnbEl7TAokVYKQo8mMWFjnykiRrslaBbydXfTGU0RTIoUEW0c37joCLk/F+vvjzr
Q97KE75iqmDF5qvCfLNNhFYTOoB7V3NpFPqY0+KlIZ8b1nC3gyBAIODeSPKQj9fJ
5POyyGvluq8J49mlnfxidwB4rFMLuCcbtJwUnZ551s6QT9RMEQvsyeNRw0xkOJpx
nups2CjAn9KuH8dfqzmV++WDj1HdkqaI37rVPdIbYvE5L6j57XSPMG9lSu6u/BE3
WnT6pks2GfMUuwjuhaqyDwmWWwOOMKdibShZHVygx0Ig+HcmvuOgho5sLrABW+Xq
r04Z6QLpFZ91kUBo4jbjYLwfFAapHGenfRNC2suBn+vGI+UGEC3JtZRVDNmJxoec
NiFTD0AVn6TECLvQ9bQ1u3f+18bxQsdrAOUxRa4/429DaEvOpGAxEdvGXsMw/NZJ
2/H9brEgYLfGAQJTo+vlKbiIkh/Y7J3G6GSk5kD1Lf2tAIr3trPEJaHMT7w9NQYw
ZX0ddNeVK2pVfNSPhrHfSpayxPKfz3K0n8xWIfJA7/Z6xylnnm3WAvE7ZERjdC1i
3laOLwFpQ+PNuqwJrq95cwSFBfmKGiBecg+Ded6oyTPl3tqVTWtx7ePZ9QNBRyzJ
hbiLawADxZYecEcFzB2ijoYMS9VAY97oWyafSjrY9+EyO66bIoZqN9LXEzzYsbj7
et3nIQIu3o3KaJGRkK9pSpwKmR8mb7xZQHMpRg4KDdEVu6Mabc4vPID1JVhOr6vG
4lFzbQthY2yQZ1AdG9CJXTHKeTRMQD89Lw0i3eLg29BPjapB93+WYY8DPMWNGxHK
62zFGEU8mVg6GvWOtfxRJ2fsRY/R/alXIa8inpCqilBpYl5SoBlouRJ/KxAFSsvh
1Mz5DKK1GtJjsOlfeHZgR7jV8nTP9YZCVGGKZEc8W5gV+DPqyw5p03P2p+07KWtU
0637Wdxscc3/n3Dt8Aa+NBuu8PQ/T6pkmyMYxVR9suTrKvqAYO2CgDZVtrXk5UBh
JzZXa9enJgUwKvvF/KYiUPTWtm99S/TuCSs2RziGZXv4xpN8VvEQd+Hn/iJYU0hx
kJs5Urh3TX9QyO1419VWdIBw2bdooN4B9fCujxxEy8D86N4Q9MdTJcZ2auSNARNP
V0bWgUl9mS0HonUTPzLlZWcG4MBl7OGcVgRcNCNqtQTTZzCsoa87lK/VBVTF4s7V
czM8mZnOYJYO0PSdy08afw9W9GUHbweJrnzvzFwoH3883WmzCNSfzzl10jVlIpEZ
r/jfRfBFKOzQZ++h0ZPHqTeBFrTMWZPaEbDc0Psie0A8j/6DsbRulF9zCKApQ8xM
MqU+qUa63y+Rf1ejMXLEU6nIgAPhVl2XXIB73G2g03ILuq/67Hmso0FEbtL97qfg
HT+68yaGKF1JO/HbRv03d8uEHQDwpAvKGZTIoA5gDsGSBBPqKn/K40rICLDABpib
X7de0K88nTvO1kBNDbQ/HQyIWIl7Wp9/KAO7n8l6mNjSk5bu/cbkC6Kobv8Vani3
HCOEQsQIGjQaKCidnGMurEoXt8bIVhUMWFeDVlRwoZzEYxzF4Mqsvvl35Nm7xv/L
GXiq3gV51bU1tW3mRIbD/PrWt69IwpX/lI1DfaouK5OFxfuc3LhpvZ45dGMp9y5V
YguFM9JomgZB66TRdA9erYkz3oWPeJHeu4jsMh927ASOcancu6bYyfwsN9eFQHpN
KRm7mr0sdU9uce7sFvHjwdKFmIJ/WVxXepd1EZozhrjORCZH7qi9yAbrWRqJlNEI
GUmTlaGivVJgE98W5YOzgqf4BkRAIoEablc07F0zZoLcaPMwB3bAgF6RQRFMg5Ot
KtMBjOzi31Rw39jyNmlro9OnrY2ORkBBkXkUUkrMLxTriBhIFgsUgob/MLnobkhk
y6aWvSddDRZwqB4SpVe1twXXefOqZrSetoqM6pqxglCSWAmmnCNw8cww0OHpZssf
+6U1+uz0wVRVr3pyFQFc+oB8p9DUApiV7HfRx9Fxg+P5TbOfaj0QTab55ecwbXTI
h7BlNrXIJBueKytO3BuJg1SWPmAzbK5OyZMqw6pCyqllbhkFZITKHUHMsnGKTgLe
YU01aRE53G5Q7Rb7REXK4YH7wAdE0R2xYyxyfII5SK1O9YQf73uMEl1qv1/jrshJ
tSHNwpSa5glCNg6imYIMBKD32WU+SpfDodCghyp+8w6Cbf55+EjqbyPG/a0GVmoX
EXeoWp56X91Jp6gciIO/HKyQAZgZG9VBgqibei6oRJCOakzl0Q8a9mZNgKEugPv4
LkiEfKMjaOd+Mq1zPiaec0ZR9MiLgtIM79uWEbrE1/A3D3qFDYwoVlWk+GPJ5jpm
ZwjYy+S0GA/22sCwqCLxuvGX7Sp1RxzfrQDVPQdDQeyBswkgeePuFOpS0vcZan03
VCESwCbYqWVa6QZyt0LGfEWFnKp50BVhNA+5slBr5uteKSVtIbrJxE6hmAm+x2GI
NdsxV0CUY6U3hor6CfohOdIvCK44yfuvoTzc+qKqKL5LlUmVltYSlJtk/DhFeNck
zUmDxMTQJRiOafGyaS91hstPtAFM/NbzDUCUrrlz698+6yveT53oXYHBOIsq8wKD
TqZ1nYl5cRwAAOGkLZ02QM1yQD+/BJNTaF50jCuiQhz9N4WNNQobR8u2MAYpT06Z
WzWREYn3P7D5ZchB2gnwdJMpUtxqsfdR3DlsHqMad3g=
`pragma protect end_protected
