// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:41:10 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
D0g1qjOLdhw3uQvJ1ThVuk+pscfKs1lFfVuQypgxVMUHBzEPzQAwZ3dmQl/oC8lq
65XyiEh7EDSvPOeOYVBrWbdROEEl2jSMZ96AsGxbj47r/Lm9sncCOfHEoDrFjSNk
DNslSLIKroAtB1rVDi9N34Oi+t84/6oDMIH5gZbeXNg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 49328)
h3HZY+EsgtyyKMeEMlr4Jaklgjq9JR1NdDJOns1pNU6n2eIQmbhBTCZvLiw66Q7Z
NchRJO3YLUNkeJCdGRg/DOJVc9CQzSohD2MZohAFau48uiUgV0wix+C1rWmlhrAA
Ni58bfD/QBImRZ0CDiyzC7xpEDTKnK+ReThc7GPyFc+FgqbL3NAdvpRGGht+d10s
QW0Mhis7MTI56qreENA5an8GGSYEF4D2w5Up4bFVK8W8qqpUDOmGGwp7edlHoKhO
ighALJBkutObApL+mZ0tm0FHQjbeJYZ1CShbo+I9JEZNICDCOgHZvgpuhiksi+9E
r2IVyiQ5lp9BSAjXI2wrEYrmxtlCoqQu3dGWokp/xYMSlSu7R1w5GnQ/xHySZLwc
//tDgdMkl3A6htg2OZ/3QBqg24yUo9QUAozqeyc2ju5gacKJjraj2WVJYXi8l/FL
KoWBlxIppwscrwWHux5O8yUSncIt6IThZ1/n9/GhQkCkzUQEy4CDBtbwc2yvvWQx
8jaJ1Iesyc4GDczthRkO4oZ/IwFyMrTDvqA3R0ggnUdjwt48U3UGV+ravDRkOBBA
3eUtqh9RWcXCgjbRpXKfvb+NjSMW77c1RdThUO1FuMFGUq4hczEqqgQwASK4xwwH
qLX2V3Lhs6NHV0kk9xKRbClxFo452XOe1f0d9cW6GonKPti9LXBrM72qkF7J0JfO
1lbr0x5dvvoOrIpdTWoQHQqpJkaYWYA1ZnmZnDIMGSqJ46lx3qJLt6Kk4LJMfCcL
VMZJIOqTfBbKeNUyPZQlSrIEM1xv72vUHV/3yFGgYVoaAS9Fcokw/XRQR2qeOGj1
RptEyKNSDAvJiq2bGaAH2Iel0Ilb6rBQzGVDFPHpZzv2IC207VXlZUxNQypSKCkr
GzbXEAgiCREsVrQ3qg1wGcFprc+0N8kb/+tWKXZ6J3Hcu5pMdAhojvnkkb6kL3IS
ckA/oUnbY8fdQeIy99wtWKsJmOBq5be9hSP8oTY1AERT9gjOfacowcAL5Vq6w2UM
KApwyNOMgmqUG2N2K8umq1HKy6D07IBlVV+12XWpGEslAGimNqmKPPOpdyncN0mi
j4MY4qKevvgyIaETvhjpOmUaxvXRL6j8LFj/GTdDkyDf1nX7RY3kP7xlLk8Lb9+Y
1413CQYHbtDHPrGAvactSLpw5+jhYbjpcSFi67bfPWg2lUo3R+04N1jUJgQUpMmF
GFsPXIqCfjiGvUyNnD/rhsThoh9WYp9ztR2mjuylnbLgt2ik8O5Zbo/5358B2STd
0ISKli8rJaMfwTEj500SUxWbAB2t0Kjh6jIWaWUhstmhvnCsQLUCaub8FaJ/4241
8KtxgxOXppwCYRLl6jL3vHGN9Bemz2nuz1+Tq5BCZMHH4+2IymUSW/N3YHhUFphU
ui/5Ea8DgKYcUXcITHxAbs7o7WXw7SzLzsxX1bVXXAsfRgUO0e0nQd3+lrxSgzmx
aOhmrGSxNSRbPZhMDm2VEYldhc+1xRbWWpQItnL5761dLW2PbCCClfWIUweTvzNi
wdyHmOsscBObwC6i15ThFFeCK7Mt2NrG/bvKpX/2R13Ab0JArSB3hWXvQi7PXeGI
i3vlx5FJMwAeRUYqEhiJgac7lprFCOPdsKY21H6U9rZmAIE8oN+/tqwHQDSE1W4F
A8L0OYzx4262xQM6bpdzhiCrmjBYzB2cS2OsT+xmHIx4IvcSH/2eux7dxjpiSzcy
uq+PVZjM6bxd2r6LjvI1e/wTZcCRbENCw6qDnh2bsFgwAbNd4v0YlROg2vFFe26n
PY2bNooaDfXlDoSFPS3PblOkbDtmFjXyvksLHQH2eoWHU8cHDgIhni/tk6II+5SU
59th/aipk8rdZzynchO9hifjFlG99mpa+P2A6wrn7t4VsNhx1I7pACUKowYBh2tB
iHtrk2LhCr/4adpaiZQYCaHo29xnUZkG8WnukSP0bQ9JDLTl09tdaN4Oq7+VOvt3
VkpZPqFuk5kCVzJKxWg7DW/x/U12IY18iY7hvvpiLRmTvF+eKXANUObG7VjY2q2P
MHon1xwjVdVFjWQj+T3+o69D1Izsic+eZQvjkO3AQR8ugwIeZnH0h8ucr434+GKW
5QLa6Kk5DAqkE0flkIixGlXDXRZqa1luXg3tOKQWoih72HTxy+VT97ycz9gt3dr5
MjW45g47m1Jmtni7htG4n3gpFdUCKrREYzS7lJUbzN5Pxi9Uq+K4VKStSZHEHyQC
7eAMr12vz0LOZ+1PdeFwAGMj5YYVnS41YB3JVUUy2IsDXLIDSePJuXq47DV/EAmr
R7ochbZbGCCz+8w72AzU426NS3qfdnJC8kCeif5LwAMYIjXJ0Hm96mjjPT0Tk9HQ
KA8qsvNLeVaSXC0Ab6Hxqm/fp5FBhsUFo83eo4WkyaCYRLA3boVEj2bFMAFh4/JF
l3KI0cRudE/8uymQm3Xcb0gr3c9oLtmJ0L+SvnJ+4S8fl91VXMlRa+B6VvkHdkyU
40/pmmKLPVZ3qe2JTskTEdW64/WS96rCTbgoC556t6DlhLmyCn07po8U4KLbQMmK
Dmv/cS85vPuIU5vQIeLM872dYXbp0LsTyf8JMszI8AQmffRd9viG/uP3cHGuTCRw
9FOt8hkRtYMCnKTn1Uw+hGEgQnSCVGho73b8DNO4ZC/Z3hf6i9auyeBWHQS5CMwo
Maupt1LeUceomRterULjwPBv3JfskZiulrdAUYWiD9w8VlFSsQ8lobg3niArT6sn
mu6+1QcKL8zlS8IL2rvZ/xv+g3/UIWKMVcpAjVrcUY+r9ZS6yd6deEiRFV7pXv5s
zVmKocMHZF8Sc/Cw0IOItgPJTjzrpoJKfuqOnUUgonirN3IyHaCbtHleEWFw/A7h
JpzkmkNnHB1ZTMxdqgGO6EKFKkOvQ0sAAOf/Iw+h7vOV3Mae+nq+CZjGeMu+7uDz
PE6EQv1rdrZLGmVFaiPl1exqE3QxBpypUysLLG3tK/WWgctDc4/duVuxWhp2m+Cw
oVkUXtDT7dPKYQdwe2a4cRjmYU6/soH9EeY3SnYUpDECQfae1jsjbKZRfePwPi/g
IELaRAQT/Rn+3kpGEDn8ZFHiV8L/W1BgKvfK+LzVWb7UodG9PClOk1odlv0E+hHk
1mVfGmYT9nuk3CWI/tEVWCRBjTaKVkepyLTZoaKULz1YSQSa1Q7NtdxTwe0kZSAc
gEjrf68iUqbRQd4LBTUNqKebWQCq9WyCyH1UxSigplRMkt3lu8JBjaLqJs+yMSbr
G//OxvGL2xvXeQKll/1qkfFi0PM3YM5ed/49+4YP5sD5Z7OHQDYmpvOFi5WRn2wE
HoKtud3LqY587azeMzhpAE7ffZso06TFmhcHna9/dJ878e6Cjso1K/i34hS5VQIJ
+S9xYWyhfaGIQ3+KiC3HoeQuYfpT06CZ38VU+BU61ZTWq4h5bwaJUSB/9Ousr2WZ
s4B/HAfNiMlLdrys1P/qTtpQcHgFqxXNLQ2MdSO1lLZ8dYi3GJydMLIG1Ow9B7Fp
xpWpGCha0ghk4fScmmHuKnQFCvSIIjLJoc1GH2YsP3/BqKYnjT5sfrMd2EvzV450
bJrN8FFyZeS+ILxptoCSiktLi2z+U7qUvlsqZUvKkv8hHv5na9eqctGLQGqGI+wZ
/D14nPZo5zxbt7kXCYuyhUxqp2ZHNMbL4QzFkA1c0gTGLTqHT5jcWW5otbgWqp3u
oPUQ/iHfBrAgI/GIFbFFcS/gvGFhr/CBpgPTAHk+nQI59Uaf8R/PeHYcwfssvaWQ
SmvOVgQprmRbphkhjTn/a4sT2AgebRl6JKmU1/PBS0GVSA361V0v1FdgCfPthBjl
DGWKEmWmDFjXIiYRRKAJAHeSIXZkmY5uoS+veI91TycCH5kNGcsj5nW7SXCFxr/w
BvITGRP3gmn4x1Fk2//YhNPdrNPUfahKxOqSRrm4tyQHAYHLrK/95FM8sYFc3ToP
/yoXR6hr1M/78NyvkvmKpcGF65iA1O+h5+o6EYyogMkFKtMk3RQQQdUG0OnsFnDV
R9hlw8jOpflb1efroQDlN/ftopRHX2eBCg4AuoitFozspx+AwrcFM/o6M/mP52lr
yz9+dmBQ2JDA6biR4Y9t6h+HhMLJQh6R+Nrs+Fb5zgfl6VZ76Ir0l14Q7AhbAP+9
Pz8GtTvPr7mxcL6pE75uVmLPIYLu2ofucflNVREWfTs3F9Jy0K/O5U2GdDy+y354
QiubQOwTBN8xkylVdm55U2mpGhSrcTtw20CxIIwYtF+CFLxqunRAiU2KkRIEQxST
Tphkv2ArexcNIbbpNSAwH3gONU5+Ri23xkG1Qotm3xnvFr9QeMXQcLaFCGwwABxf
YHCHqDTd5Zj93qppBFRyhG8gf+XTQBDR2XLUVBStoRMsPGd+OBGCg7GT17PHJrJy
4ELfZyqVpISALOZBrayI460H/F/WrrJhZzCmCYVsxVRpQwH92xqz3wWgmVK91TmL
5/VX5YAjbv9UOxr9lrgRUfuPyerTcfMi6csnpvqTdcxJnMMLsA080mVllzpVIdEo
VZWuJcffZbA0VfI5snyXPwU0ACzn9okVBSnFXqSJbaI1GIZgCSHngq+i87CDcFxo
vUeaJO11hSUNQf1CQbGJwURxkWEEuEEwDUbapF8P6sFZw8ZcyBrb5Weq/3t7ST/6
mWelXe7ABV3q0xcX+NN0AZLSAm9Z5FSkUNY8ovg24U9jx7kHx47q0a1GlH1C4ci5
Wod4trS2exQUGv6BBv2QgJasy6yTth4nklcIPFOqxrX+HOV9w9CCAJ+c+16mQ+mb
pFaMHZWSB4kVWCIIX/WoBwJjDyMnvxuo4spdw48q+fCTf+81i4dBb+WyZK6CcMDU
S6LFYGWidBBMojiYw+BlXwr8FGLCldlS8OAG+VoZtGBWXltW3OhkwgbPEHcP60XM
VNI5PIt80YY0ZZic7siXU8veHQs0ErQJs75J08M1rS1QXiC41noH3fgpkfi3TTJZ
YH5jgXIPhclodjRJLt+QYl07BJ8pGoniXYsvfM9ldkK0ZtSj3QXF/BHcqKksMEDj
kGFiRSKvwajbWikfPY3ww1eN+9BUXG7qY2w+NlDg7eWZoUSvyJ4mg3BLFyaI4tKL
6xyimBbGKNinuCSgG3pt143h4Q5ILpBZgG9iI/5AfvDRw4zcc+E0PmbKecJl4t7A
4jX9tiKKgIcMCebu/hoCHJOnUCJaVL3FVmhc5Tb+B5ikLkt92hP0suiWkPdIVk6g
5BOL6C7OCqElN/2peX/dNb2m1el3C/WsHqI7jQ68HVu15v4+4JPe+EhlmAtoIVe7
XVoNSNuLSSrgTXX3MeGfNnc0vcorExLVsHJ5oEebk66uC/eC7io9ozd75pTAPGuu
A5jCOe0R7QXQeTDZmrhSEYVc0MbVBuIeMoLhyZKa6GJAnxGcKLwBDrm0aeDVV7E1
i+8DUyBT7kkMfJ7XVnLkdwtV6/1I5dAjyAJ6vwFIzyWPhtpQg3AdHrIXd/HcoV7Y
zmlmMR1nlS00aH6cGnM2Q7sCEcQyuc3qTuZ8m3yD+CSeS6x6aQczwghBL0872eVD
Dx/HDlXSrSHJ8GTqcHxp+2j0MEvtoZnF7kaikyUZSK+1cdjrDQzXG8eFjK1b7e0R
B88tYvY47CS9nm6YFvWlDrVLL2c2MEGx5mBWwOiqJa1CT8pVmERWud/fhnD62ymq
tEthW2YtpC86RS1VzPlcl1dF4a0B9XJbYVod34AOlEjpmNX6yMGdWisycaVxe27H
FXvVf6mgkiV6UfXcBtud6L2vRl5m4ZitvqtT3pzzRdr5Y7Nwjfn3NI7OYOeaQXjZ
AdJFEJx4/aogx947xCbbDMMs8zuwLS/HfLoRF4DpK8MB6eMvG2MGakpovEWWs7h2
0kSDO3j+5Kndc0TEr8VVzwdfqHy5t2cTWIPX1LdF6xPUzZFcwQNS4iC7afJYdx8q
K5ptUd2hOlOqnTunndzO+ZKAuvJY2l6ilPlDftonjgIsOVdlTGz3yJcyGgLvMDvY
0WrIsmGO2bHLWsZ/jkEZKdXgCRSwQfUPo3zaLAtl8fslX9zscrocNI3HQOIfTWxO
Mw2Hhp+OZrhEpC78bRW1RebUn5brzeTzoRfhGphpkBZDu6dWWRj0fkIRc0rh5Kxv
AyBtbZHLThmdkpMI1GsLa6EQL/EujQomXeXv+gLjcK/2iyVl8d/G3eyhTRpIVIqY
eVf+PxKUkjFhlYAC+I+kQ7PEv5kIydL9kzsm2O7UW6jbJ8Q36RohMcMoPr9/tYJX
gL0fRIYPy2j3frsgVeOvcgemtmqKvrcDSue5Is7Rm9XkPjn3YXgOYjJUyj2yNWEv
TXfhTvPH8rbKgPZKxDvjRc7ZmxwA2dJihZ0IwSgS+DR0I8VZpGEBCuaWqGQN5bml
o+tRBB+wUGP5fzHaQjcev+Ieli8DKt4b9rajHf1jvSwA96mNfz4/DuHkNNk4MEje
2pdOwKmEnsQ2M9AFgMCLiTsPFyzOUzeIyyqAApDcCfBD73c0uAN55BJsZPl7ZT3f
bKpTq0MVapUpGmznIKbkBJh4Wbe8cdVYMsiW9WCjX99Tcouyzx6V4QFKuJMkX0Io
YENq4pmFQU7l+j4mL+xkw54Tf4gX4phfTBmMs7qSHlORAciNHXVuGVWtGzDmXCx3
NsA8ypAscs841BW9QwLVSHtN377rAGjHbvlUWqs2lY16+DH4S1+Py226enyTC/hg
kJmeXxHkHqhSV89bINibWEQNlXqEGfLG8a6IjQI5NnxKlWvL46TQGGoLc4BCZP4K
g8kf5T+ihal5VnfTYXXn+ewecyLiVpLH4lILi9NyrmI7duKx5RSw2JMdpNCAsdhG
a4+x5uYJ+HevNHOAsmpjYRl+vlsPJPRjjJphSyuyGb9GF2Xk50hEZl6RxISrNkYd
T0ZNEPXUWbiN0hvyH+WNdHPsoCau4MYeTUgGkPqn0SZ3tZwnU09Idab8bgcsf3Mi
+3fBEP0VsnTtWLmboCSzLcCy0948nefvqSnrlZOsBpi8ML66qX7RIpQ27Ok5R+aN
juZQV85FtEHwPIsx84DI6txyKdnj1jWQg4a6lFFQcYYaLXtuVkpHJUHxLgXqN+qm
lIkLrql1oQVMYKTdvSxa5jbxWzcYepocAppPCQE1lRVvVoDz0PjJ6GyLMyamJ9Ih
Etat5LWjJWStIUtIBlkNza/yrovlgpYfqgWZPHYmlM3zIeEoFTwMgj5IYb8aMo+n
XhVdqKLFoClz3udh0sQWFnEIUdRlXKRLfyhUOOKHrNS/yoHZ6aYn6r8BY5bZm1of
qjuPFC55Kd0fplvgD3Bj6Nmyj7ptNHaTlQIJ9lB99cng0VlcKbd/TbhrJ0l9fv62
RuqLI6ZigJofeBbQDb24wt+RHlyFRVv1HegE9atZ+jfnrXCM09+8QWrQZRrA7nB1
AvQ0vjOfusWLm6Rudeg1PRS1hv1nP58mbH4lZLwAk/N+Y6/uDVK9bUjcYkZC8gdr
OPZaxNItNJsIU+Vbvm3b0BguT44SMAMwja2jnaC4UNIG3Uo16PftH9UwiYSdZUfo
4weHTy0UBTgxmESaohii0yy9Iknq7VCOp3Beo7L2FxF6U8nzk2NhsR98eWI7qzvm
itSL1ACGJzHZfCwpXHMm1mYGavobX77l2ZBHYx9XIamfVyvdLIAiVuchzH6bUSvg
VvUCkJBMbr2C0IM4V/19xe8bi7cIsSFLs82Rj7JlrRAh8hynxitDk+yzbPSyqG1y
rVuIEVJWMihtH8eCX9n6COkUN2TmxE6nSsFFf9clrf+NX3fO1L6QmVKMcTJn48rC
g+8XUWBKAzw0udGgoFERtUJw4THnE3i3gDqN8g7Y6h7Am0VcRcVN0yOk39lpBqge
ZpLNz4nWWexMTuhcvu5bcNsqhWSezjyL/Uidhu+gM7y84jGgAjZTs8fRag7mEfCM
QfaxdOO8KPAGmfcUeugeHe9VVR4PG9JmSFfDxajrfHXwBWN60dG33MMArbjhb+vW
4tK+UzgylKU+jvl6DipWxPJzzPOwTy2OdODrCy8PohIwbaoMswgSayv9qaPHaVw4
TC2vM0YzIcdD4OqS3sgxin+m8B9LeOX8nqcg9uiaT6OSrGemwaSeL7mKaqzP5Zyb
p2NS506jBn/+jswbBkLxt59A4oYoB0qAV9QHUXD4Ixo6U4dXFiLb6sWRxX9+cKUS
0OKx0mez757jqE5QdBhCWtuqhSW4cSeCnV7f4X+JQGoC0vHxxjRgrSQWkPw5A101
r+rNVmkB9fEiSOf+uTgti+2AMs0K3EESeE+fYErn9QVx/VvHtvUc6geLzFr8JXEk
ImRb6faJUd0TKfeN1v4jer8QvtHdPU/9UTKEKHFSuF4Y624ZUIS7ubqJLwtqJoim
hOge3Gsr0vNd2XHW1AUbSxXeM8xTJDsJC1NamrhiQJQrN+hwG9bGuEBMxxyjT1r/
hI18fa5i0NIXB9e2YfvtnmieoDQJdi2EuKcM7CQWq7IyqAUPH63UIcl3Z7j35r7V
DCfWIOLWm4Wu5KhFNNrZVPTEHd+r3mWr1OXpk29W+K0wHSGXIj5P6vWRfLhIHLoI
52Dt5riO2Ko9JPx8adK7klQvhDQys7MaQgYv2MosvTLyQWWknivlVQWkkC16BFai
YZtria93GMV8kGaP0vPCuqJ6O4zOIqe5DWmlT5JYbnW7uv8ZxueQ0/tbP/AE3S5v
B94RK/d6sblrYphm2X08vAmbvNBZm1DREihCzj5BBDYXCXX234O213aKFj5tLzx5
oCXdqJsPS+ZWEj6pHO06fD/Zkm1Wj4Bzo7PMlWWsT8ZKnCCx3mZV3oUn+IlsKmUc
RZCJS6ZUjbIpEGeTfFMMp1K7GdATtUkXYmp4bn2wYGfHlJvfL8rJob1/wUlOIdHL
N5FKBc34eQAnEKq8q0tvTJhKWjr1ZrRY7NV/KUUwGcpd3jwp6+0sRszeLK1+s4hG
G67Dk1RMpO86nrSKV+y/lgjYQswHfMzKAZ5DdxB/2cgtVI7Asla+o6jxFQADOFrF
gXrfHBEjrzpZdgfL0IlYAbeBh4WQsZL0ipQ0n1G/Cc11B8GIamCpqnOcOCrDM+Qm
+ILgxnOUEp4u/TOq/DU3pP2vEVrL+uVjCHFJ/jGRSrVcSoNvLz/GZJYf5alVSlK3
ksYyCH6dj98+O4d9jC+3OJqjunyAi2d2+nFZBM/87gmG/7K/ljyMD8pi5oOW2Tto
4ng6X/bzyWjUgyIFhxFWigLOApH2tzy4JfS1skYBR9Z4EyA1qgQ0pKPc7/lf0xFG
RcmsqFzLYLTgWIZXYSOaxHCftL9gQpD9Ajfjtwu8fp3UOVOc9HVfcsvjB+OK/yGG
OQ4/DWL/H/RCj0a+jCi2LMYtxClhdZexVEA4fPBZXY4cW8Nhc/EGpO3cBfPjSvpt
oofxCZdp6Tft95P/lyTWFC/1lKl6ZaaTZi+lSADHFYRxNquQQDwaEUqt9hzn0Wp7
r/NrWQZCx8JpFF15UM1g76Zt8xSl6ISeD2+0i97naR5SiXNxnFXpKhMDX4ow+1aE
kSiClBBlU0KsuI2uXP4K5J2C8e2a9RKkfFuKJLEEGVESV8mclurswRERFVWqdHyd
dGDUpC3JF9YakoEehPju4ytDwi+dO+AHiZ57NDMWxvqRlBVWhYgbX6fTZ4PS2KZc
WYoa3C/yIsaePvlIKq6Nd1nmT8PiqGuJQ//aXTcBl7rwVeHEu9Z+YMgclz7A1get
CeEFv0kT0QyU/1eSUDIZ+BjxTxsO40k473WHeqxA179gzPm0egKUZbPIXHEJx6LG
P7Ft/FzoVEyysL8t5TNXis/DTpgy272b1yPLBfFSsaQs2qHk/zIUv5YDxmVQbgHS
+WpndkyAuptiuSoIVRcjvZhhYqGWakAYNpgy8iFNyFW9T/HROAE93BKwXZEEV5ra
9hxQZM3oYxQkfDJVr7hwgNrtXlAbyBPZvjbmEuMjwbQGFe43mnAc0ORcjjDpvVDe
XitHeWrtAlwiwFA5bA96pK3sMVK53/xQHO86U4/BmDVR1w+ZYhXk48/zcvjXs9YH
u4qscKjPvKDpDzcePYH0eU5+9xAbs0MwekJb5EvQJVpWxX19Qr9VGfEFuenLpBtj
nv3VfvvjandiBSLzzkN5fn93aVUJQ/3cBGt2aerRg1UURMTaiTyIuu7RJNNmEWBP
96nlvZDIxE8nk6SmPXFVmQjA5d1oIfoPHrCCmgqE/beAiydfpKmOWWYekdBsN1ip
JoQ4rpn0i7heP8xvKRXcNSkLg3DGd/prqEn7w21w88DwIWzYZ9gqnUUPSn7k5GBD
1ezgOhR3SduhRNI74kERlbIqPTaB/wKySIzyQNu3CRu9FscP2flZCtnF2to5WBTG
iPf60x+n5cI18DdvrTzdfmaUky30L4mLE4nbuIDgk7OEIy0IVgCsGuy58I60Vz//
bYm5NIMwcP6GeHBd6QA/n9YQDNBGC5v/5NpJgOXRFLS1ndzx9ORCPoXGcodoupYv
9pQSO/PLCOU9BkEE4d6rhUiTYmA7etpcYiDdVXrvaSemIHIW+NZ2uiCjvsyJs1sA
Ukklt7l9AlmIr3fFxLWwp7Ssou3D7/TCUnzBIcAvFLn2sGPliE20v+C76diqb9FG
N2nAiLJ72t34dzAIiNgw5aqS6f70EfWkgMGmP1dnIb02J6Ik1U1Wlc8rAsbps+TB
lugD1KLi6mLtQwIXm8SU5w4+D9PxVQ4Hpc8LFF1N4fJm3ZQNscLuQ8PaGA++O9j2
hq8/R6kNez7rg1ThvXuwYztFtclv3CENS9PGAaIeEnb+dHyw2dF2sN9ktIKLJryF
vnRbxnuK4oEuyKxNxCkKRBl/aDOa1Q+YH0WC6sqW3BX8OhVNbjD/k1JrtxfDNiQf
eI4ZHOTdaPI6BAJLklQEmLf1JJpFeD57Ens/X60C51ziU9+HJE7zYrwGAIRPV2Ss
//4C2QIaQG4S8Lop0QiCRMi7V/GgdySIs0iVBDPIm+M8MzZD10IRfGbPs/2eTReb
AgcbU/hIIx3QgB9Z6HdrqZRJERHCK9S6hHde52sIelq0jby3NmAIT31Od+Sc3n+7
GWdZXiYVqd5lFPqdb1lf0k8szWGkec14zk3jUhpbVNSxPkmE5IKWozBLBWxzKL/L
tL6/oxCSSQQBqpelM1zyd8bhW1r0CFrLJCHt4QWz+o2t/HEI0voDMrHtvuy/N75R
X+8TTZM6XweeCgm1RD14mwtoN6ddAXuoBt/9/GcBTfXKJpOe1q+4L+LtcMMHNBgX
gCM58uDze6l23HpCeh4QOUcS6KSEwO3JozQQFy9s5PSspCI/gBEMCqtnnOh+m7EQ
/aB4OZjploRjzYzVp4fOVVOxR8WvoLr6seGAWW1HfUOWm8pH/Ih0X4lc+PAFH6+O
uN/HWWlzL/WWvcdgKhcRJdeQffHHrBXxZep2Qhu6lG6vmpL+ay4DqtzTBfOwv8fm
OwOHBLO1OPhAO6lXDqc4+lQsU2ZnXLmlGD4xOLT7JTsntafsAL2E13yZwoIVf+TO
h5HMwDW4S5Mp7gO48DOJQvq1dl6Hwh7ZjSKu1obSkYDwexu0jNoGuy5F9KpgtQYp
qmISaf6hkMfI7PLvBkuwq+KS3NthP3JC3lCV6EBePSvRu3iFjrMiM1mqk5kxr29I
a1acT2jZIB2Q0vw2r/+R5Re+NzGAkpFy6VH4tskdupqrgvUo5ZxT9rZFJdXIOchD
tpr5VHqtZ9bzF4BO26qSooRdqn9TIowcNniGEvsrfXIDxy5Kak9g0Dm3YBho+OxB
4223sVyiPwmeHyR/pBhokgbp8Au2nqVbwBkQdjkpqbleUFj0GzgMA1gFE5PkOCS2
cOhlsYlPDnbQ6gThmZv6ydfjBcutqY2nYUFwoHFL0/ZFgXHvRYEEH/l10gdvEnm2
GSBLViGVGEWAosASxGtGWz3jCXy5nKei7PpLXml+PNNwDarVBWzSYqwWEq63lUQ9
CXzWxlT4+gCSDclgG8ByYH0sDeqQKNzFizUEeq3GvCLMGVSt5TAti/6kjWqA6LZy
sU3Iw23LkkwEEsgBHl+BM7/HEZ/5POJ42aMV0QaZPE3eREG+vDsfBztuT4n7zjGK
cthTNUxoR69OaeTnsOL2Jhn5rFRDQ/VwZmyb89beOvS2YZbnms0B7wErljionwQP
hedfHWBmUqWFZk7nAsaqB2Kc2ggydY8BtayYK4egqRl/d1UPcZiUGkaLuJZcjk6v
S4DXnsffTHBOOYegco8Fo4sNMFqKaqN6Rxoqld101dwtfvHjhHvlIO8WrVYDdRlP
AXnRQaii2lZShK+XDj5ErxCUmr1fwC5duUjRMxHI8WozhRx2IiSf60yZd6238NnF
EfBJca8Qf7Y9mqPYakdcLRPDEPcW6vooCXCNwfS4f4Q9zx08Xz+VkfGXDc07vzur
94Rn+9yK1XGizqGO0Ok5EshfujTBr/EPPmoGTbjsUo8HnmpbMAjrJgmxw/wJpgJZ
bkw5rGLTS36MrpEdNA48WLtzJc7oa5FoDxgt5fxdNLmwnQELQrqeRFuEfSLGmQJo
3ACfUi1m9uGvieOH4W7Czr6599DS2PzP8ROlpTp92aRCLrF3bg3eRv5Lcac0ycaO
MTiSJ0L2DjSkYI/Qrcw22QYcejGqPaqyLvtZG7RedHzDrwKvG5ZWL25KKJOi/DRu
+jD1KFg2U6nEnq4vjzAWZLJHBuCD06fTs4jJ0JssVs/m06Tj9fwnvYqjXJX03YHL
wg04YItO5z/1/ZBt7LBoJZ6P8NeeVntbgakQNDKlAtPAH2rlSCgpexEu+sexTSuE
tzYKV1Yl9orBx2tx3nKUKN72e5c8swc0oJukLGSgixoDShXpWxKFBqXwq5pHEhKw
XHjqJ/9V2nqTXU4QN8OJtj5FNyXuJnvEN/Zygkr9ZbIpi7yiRt2Z2hjKtLjjyYGG
oPvr2tEYm733WLayZYJmnFCVJ++77l3X/mRxqRoDxUJlwpEc82XBG3QP1CoaeRTX
HCgdhrUc/zBFtFJiFyTmVJ1X91V8OtlTO7tefsizZ198ytHpo3aJ7LAzDLj6yvlm
+PFiRifV2h06BIO3oQ4ockcrD8izGD7MVz1Uy4yCy0RR/6YdT195ergUgV9Ritt+
XkZpWCxbYdfbDAfU+KI3qkGcAzErTsKBqQFLJm7nlJJXbrgmqMDia6u8qJY5s9bD
MI1JMFoKwj/ucyTrBOcG44QruNILs9pbNdIMk4PgBd0PDdcy2dl8lRUjRAMQWclc
CDS1BJ5DRfuAEYwQcS2tl5SeR/nMm3/S3SU7KXk8oNi0WYkLyqSONEjs/3tj73AF
uCDEDHLVcPuPtJoEYEHTp36+UA3fZz8NGtuaMllg+vdmABxS3h7W0a0t1MOrQIOO
kZ9d+HBt3VnlXeJwokxV0Or+x9XEQV/vrSjXNu06GvbakutNhjUpBqfUK6DRlelf
xi2E/9nHyLZVmBdGqg8nigHcRjtB+O+3aSr2vBRXWfbQ7TyNIBPp+n7X/F1otKIX
7fmssTdLSwVjhPV5b/lttuyrdbM6tqnq5oX16AIVxIUzOk4aTIrV84fT27BIBsXv
7dECKf4Y3J8UdfmxFwXP15qY8HdJlFVtONq/35LSs4li0nMJQgTNmu1yj3hc0ia2
pdqazyd4Jm14/55m2QColaKsVjtWjUvHMUDmCd/e0soGo6nTfPrYGjs8895UKWjZ
jsWd0ON9NJt1LG2UZncngtK4iLlotW9aGPEY7HhHAjwIwLAq5cF1jx/ZqlsQkszb
iJpqFTtVeOJkZZ5o5htXzOavJuRrufIuGD/rYnrVwir41e7ccCz5z/CtufVfv0kp
dJU/r5Eo7qpNt29hFdUekABZK43tCve/Q6fkCnjAm/FkL0Fj5VVa09kxFXHzBYmo
Z/fhcDk2J2gtQVwanxR+6abypHEL0QOUcNYBr0arYk/tl/Y2iiYsIBd4IIbxy7io
ZKMjMG8tu/OTyXz5Q+7OQcnXqZhusShOF1+S2fNkaGWHugtM/nlBGqmtrk3+5dNU
oOMjNQ22HC1h/4BtFl0KsxfyI+l8E4fhaSHJuPnty0J7fdSlrmMoG72ogPu6TIrQ
0LTY98F2ky7wLMna3n+2FDPScqI9CCtZrG1NWI1H4FIUKiz3YovqtX8SeotFjL4N
XgWGE+5WEoZWM01z3m5YY7U5Bt42uHL2KZPM8D6ycl8VrZ+qvR01h4K7dzO/FQUk
EfDsuJrBZnLhUFrAMRin0lRFChGI3cfCUSI88MdyKhXTBTTLS1xCtkdM2hmrhKng
QoTQXHUSXNAvy9X/6tcvG+F5oiftrU/ryFXKmD9BynxGdnyHd1A6N/TJ/LmIr4GT
o5mP/BQ9DeBFXQkHQngxnAAp1hAktMkumCq1dinR4q4+70Rod0f6i0Lgk2UyLOZN
4HjewyMg26wErds208o8iuztHvcAfx8p7C+cnW65r1GEylLcPsBup3et9TM+O54E
4UdX3iO6kx5wgGSEAW4d/0pHMXSmGw17JVZvwiRGgkdmqPYvJ60xn9f58CoPU0mc
sS1q1rcM1ZdWMIlu27rO54ICMzeBE4QNNbCp6P0hREf/8C7fqDxFIe+dA5QaZqDd
OSiQUlQo5qUxcZwL22GTIL3BeVfd0x8PUfqJdgauEhKC8yfJecdVVUj8LRqfiplo
86rHqXjYMRjOOsxvJ1ofGUuo8u6E0ITxzoMae1QHiiexLVGzMcYuaHRorLFVipZz
SvjAlrepCGRHgdpxj/E5FIiG0LqN109O7X14dHht8nPskwVtyUlUFEeB95qqfK4/
LDsQk8/tNqrYZ0th3o/IvCz6Bszzh13Q0b/rZOrRSq+foqs6RXFNfRZy/H3gb+jJ
ZzhkMlizNnKGnd3a0AL4MeYtMOxMPdeOzgLoUX/K7gBUIWHh0+SASx4sLA72oS+d
NlFB5B2UxlHtqgvJBDkiioFMRX/D8ms3vviBX15I2gZzpCWl0MgyIX6JVhVOl5e7
6bcE/Qw0jU3InpBSxWj6w5H3Ck/8x0TRMruBAFal803Ib1wsk3ZQ3IbxGd4QpB+0
ZOQhZlm2EeHeUCdKBRNTJmyoYs+MSrkrQ6JVqSsjOfAxG4iEtgnsXYqFaUkqa4vX
8ADWNrLZtEfZwYJtyRTDIBZmdI8HEkuwFt3FCFOl+hiN63BXwAt7KvbHXaSkQnYr
okz7ip5hVbECwDphttatkGTwHl1w01ZK19WUruZbNFUsdbfS0sr1UEnDzbEA8biE
3joPI4xntXEi3T56nK/vY7Nvt7ehwv3t+7Yu9fxNyDMUy8PYZWj1IXKn2SrPKZqb
p4I6/5KkxaJNhBCi5pCT5lOcLdZai9ZUS5qOVX9hkAzBQGPTvBScjUXZgIc/Dvw3
b/teu6HxFfQ3uWUmJMofPNd541B0MaOTn+QIiwIm+NrQxzvmjhsK5GWN/CKW58vB
053odZC6+H17pkx9ujI5DUMDaxX2DW1+VHYo8QIE1K1hanTCwyu6oOMSs2YrSkBU
dm8Pau2OboMIXHgkJgRYqM+lO0F/5LYqseZceNN1926vKGZskMZrrzIJKnGZnJGa
PfHHPT6mmK85FMo5tMlZhpa6jf1o+D1KBqByN1FR4nvPB9MQnT+9FGDRZVvffsW0
q5CmUWUXdo/XUTc4jnU8I1zbMNpvqpBa+u4W3vaAQewDe9zDWyLUIqFx7Od3OxCh
jFENFfvQJYQLZfbEPBgdlcTCrhl+cXSh1JSoN5FFKtpAX6+YjTl2O1cGfaUWdumY
qFN2JjwepKz4f2usfsBawtqpZ5hbyLRHISAV7gNaDfe+yhqjCEzF0hNMv+CeMg9c
4IcWmv8PedWLfczVDKD5KwgaRBgB0E3I7CTxMVC0seJeWCxIbeI/fhpmlg6dlE9G
OM/Pz2ipYNph81900NCldHlIIrm2abflc+Ajq+bQRt6EMRjRtNwjIvire9CC9SOf
NqxLf07i8loaHbHRcaVmIvnxwWxsBU8P8Rr1MZ+vUkV7wJ2ec1/Oo9JQcY0neOaL
wZXk61klE7fV63/ufoa8qV6wJHrHx4htKCPqD7558ZX1IcJzWNOed9uggj16Bmu8
UfLbA/A+/RmwFDpU6e0mOyvJsvh2AyvFpiN0A2+ipsXIrRBbqJwKOQVlnmmqgLKa
rFjLJk6XHtDtht4qYmD2ufqBB6Kp64g5KHAjUkjLfiGU5f23Kp4h/Pd2amCV7Nic
3UUymgP94p/xz5OBW8rRmiOLwg3jBmejmN5gPwPSvHSpZFUN5sL5mhYYiMPGRQYZ
gQCuW4HmPIGGo7F2S4f9ZYbyqavbDEv8cu3HrJ3Gs7dynSB84E8Z84Mjkg4i7wjg
QOclUz878zgfwT6SiTHn8vhupLGPLQxYO+pgzxaxqA87Ng8TqTja4I9LnsMUbNPa
Ps8FY2oWUpBb6rVoK+lyEdlkpPAggRiaXtvssEyNA0t8oqJExonruc2fFopSQQZl
KPSLwtPAqc/AOGYbODtbo5YdU6REVwOF1EHDITNV6u0hvv+DeEElPkuhgdYfVoAA
r4Ns3BXlPWME5Z5e2tqoTKx7/RGqQ666ijLXMhmwp8XxARSbY0FHG+w6z8GAc6S9
VGm5f1CfP5UYuKqIJ2+qrgwI38eK+vBKEQlEYsDQ5md5rfs3a7EpLiR1WfVUktTI
mrufQuH72hPcQsJaqGe5Fn0P3v5tMMkk9Qvq6fxK4CS11ztxQNzqDK22rxUsX2nU
Tm/w1u9mbmzdVxDxIssc82pA1cBw3sE61QGy6g2ddlbpm/uBM6xTihiAZ/fIr9ZM
ddrEfw2KbkC04DFfLmAh//mgLwTvrO0yKmpVGkvNNVLM+YXb3LU5jBzqSLpR3yn8
iIxFnK4iqycNDg4KKV/oYQbb5zFDaduGP/mxohppfODyLc/vo1A6TpVUhm+hoEX/
2waYWPXWZTFpheVL59kJmDbtvMMsi2HDUANIGmvKiPdKkAOeUXy9Y1dwzBZSiN2Y
fYkpNnMX92n4IiNJGR5yZ2OpQX2Mq4ImQuD6ri87S9S5gDkxr6ZXVNcHHKgg34Lp
1zjqm1bIi8DkmejW+GVHL6edLqJcUcXji5hIL0sYQbwnKblAXOfzVaB0ZqftPOKq
mUkjKJUQ84dI2mJlD3/AA9Zpebe2GZIyW3UdFXYsHuTWvVanXmVkhRh+B8zW5TGI
HBvmx8tinqwe9fPjB8qGvzzsuCIe6T/gXd6IEryIQpWthMiT9EmS987CZgVlFRnK
alwOhRz47bvvt4aycQlfAHMlFRp72UsYTkCQuw9PcYBeBQbDopXKgWKRt5tQ04lE
9rBTUfqwzI5SyMrh1iAwT21BYumFQHX2VlSwQvfF1h4BEWt2avg69hvzvgChW8QR
Ukr676pRJuJS7KR/IB0W3pmxIX+Gzn6w1UI++GduPS8JiPiR3TdwO+loi8k8I40a
lNxPrO071f1S3NSHGRU+jM5ub/IrzpRy14J/OeFgdMwBR8Lr6I1jxVZeHhV70qB1
wK6AfEWUVVhikzZiMEgRa/apeOeUmIUcnUrvDcwOG1TBZTNeut1uaoJTzP9crBRi
kBKYnDUErrXUSoFMlEcdgDB7gOiVy7FBN5d7aclEm/BiWasovN2mXHS4flcRxzel
sETRGLX2zYfahzrtcaHGed72QLytscrwD5zU8IT3fGoI5QNb0BHLAlNlI7OlLmy+
bgeutbpvTW18XmnuBFtJIYZPgqs+UUQoARo3+NAN5mIVewNNEUkb4jdg0vl0Moax
271qCUW+vaZg4MMPRJopZFzUhfIdI8ClU4mtTT0QeRJXjmehEQokX/eTCf1G4GZt
8rqAHZJfe51EJi1UJ0Kx6GWbIzBlAB5WxiHwKfznUCuGlUbqNPKaJQrtcOgd8mpT
ibqaT1dYGacSwuLQzjq4E4OpgAcoxNt05IaXZMxoNa2J7kt/DCNBJ64lpkjiE4vM
Ilt2qs/NLt0t7vxyqhHpHyXqXJvieHBWxzK+dV+M8VKUOrtjCN6KjNw75YhiN7Pt
9/lKQD1LA5UWCuEp/htya1/2kzhiVDIu0icMLcYu5kh0byCxnDj6Y2EnXtXizgON
FqHuthcg0DZuq2Qm7k0Hp+hJZY34jnpFkbgWSrL08A3W9hU+XBji+HFv4JZ/KqZo
mCO8LvnQZqhDx3d/HuI5617qGrwzO9RdMj/ML+1Rf54ZGZUG3caS/kysCxnUc5rA
hqhy8+U1APsoBRKoUJbovpLMrqBoK6DRBNfA3DeE/JoBmF+dd2brKhOuSE4U6sRX
3BagAY5xPvKtO09ww6Icqt8SLzRo9OXeX1S0BxJ9Ekr8zaCsiPpdSJEcCMN3QhUp
ZjQyFhcNSfoZPgi4cOzk0CXAhGAYXaSHj1/nKxODPfLHThB/hbRE08/emrsINTxJ
1bcFKKIGro30XMuQEcIsRKlR0bWfnKw38nh7d9+J6gnQQGD2ip3VQNi+1+MKqRuu
loeG69ohEHtm2aUJOeR1GnQJu7mKgm88Z/ErNgF9tibE0eUBxEX9B5ZIU6z3p4b4
b0uHZlxR+3BDO8YTm8iuu5f3lE/aQ+C8fOUeop08jM/Cxadcw6/U3ghbU2F+QUPP
N4xiiD0mLHJASZL0Js9AL+BARWPbwAwEu1jLM6HbSZqreTdKmIgtq7RVMjEhhrj8
GleRJZZYPCv/IV4r7zq2Wv4snHKblQ8cyOYnGj3JCANcvDWK0/ITSIpcjOEYdDCE
cOhlRcWXfNyf8VKALfYjeuqX2ntAzQcyuqOoPXNgfM8PFQRz2EIUxxru18tav77/
OqTOAFD+Q0CWj4jYpdsrXNJTrxZ4XEhRITGvDaQtL0oMkTzcLy/rT03555MmeF9W
hJT7xZ9KtA5QKSQ1GmcEiJkP0TPPATEIQ6pxoZU/fSSkZy3R4fUxmiZeYIzMPjVO
+06rb3juc83ac4wKl36dHlO1jEB88O6T3i5yzWHfm9oVN+vYMvjGKgs7FrHAzx/u
D8AVJt7ObVJRHMiP0/rGOr1q0xfBX+//wD5mby8jJm1K1ayA0fLCyqeIuN+lWKiy
i93RQ2/qd7uzgd1Qk/PxqdFcSlXHLC6yWFFlXofyfwwou7PnGyq8rBpH58+xtYPJ
PsE4u0/ZwHUKTMC0XvCU1VYTEsxSqEtZ2b48uvsFlX6AZTTzn7UujAwbSFrLLEEt
4F6hdsrfmubyd6VJQpL0lQJ9v2Oo/jeL2hSOFk8SHvagtn3Rb6jfvSsTKVKvUcAU
58FVpvRB87WOddu8iJApGtBYXD17x2dU+4e6WjAcpDnXxFjKaIbUFZSASKEtemNp
/BQ2sSY9eLuZtSdxc4Dqo+6TJV59fidcDOsi4idgRLttyiC+/5fRnoOAwdtoO2UJ
Xq5EZ5XpuvzXrmYzbayNP0vDxMoOT99C+PMFQIJpp0xJhrY4fPfaCwN52Rns/Gfm
FOvrqKSy63ET7AjkfT5t9SABnM6qiIVPN9HWLdEYAcE13PDmXGacGXzPVHVIjAXl
i4s26112Ghxp/Sxm3LuQ3hc0r7gZoeKwauinVSjvinWL5Y/er2k0VHbXckvxa2jF
yVsKqyk2Ad/njIbEtH9dD7OaOUnCphpUuVGWlHNnWVkyARg2yo71bM7kjqskX3DO
ugnNty3+LjNoCj3t8De1COhmRpo105DV91yTzyZy8pb1xbmQ1rw0iTeRGwGI6o2M
4paW1YFQD5dRLusOSmWolH04SsigR31w9M/TsPa0YByVK3/AIQ1EHXXbZFX/MpD4
xnkdqe/8oK7C4E+tuN4XjQamXBqO/rMPpkp8/VifPwB3Ucc4hVt3ng1fgG9QeNsI
vfbQtteF93cZn94BCBoZVjGVpIQKw2J8gqMqg8x4rSJMV66PDy3MOAv/Ffb0QbjN
17rrmjG90xh33ftoMx5QQHXNcKNSQKTfAljcAAT4bcygphPo/K3eUl/A2cMUN3vw
wXgcDrVIQQGH5KYOhsqCahx0wikmjqCK2hWQt8ms5h2/qcPA9qdMAaPWZiMFCIEM
6tOSON1hIvK4HwmVC0MOTxISMgAq7y7jNaNxpsTedxXv26hlHdn1LRe0DCV58bAV
iCvlb0ofg+obKpu4ZqmHjDKUXE5z2sNR0SMy2stkLy8sreET/VU+9Jv5AN7hm7AJ
Ryiu+ZC6sj8mDIqoqDZET4ICQTSj4oOHZd+TakJB6onf/3xU+O32hUivMXGf92Zo
d7aqvL+aFq3npH1+BDk2q2srFJbWXuRYsrJpYta6norvUW5XvgsQUdIe/DvdK/Mq
I1/2rrrz3Oyz79wuP9HoVvex6xHAhhtUyOV2uKUl66S1eSGd7PwKSYlxLWu5ss9l
K4o3bCO1Y7OAHiPJj4LC5u4GV0rxiDV5N0aFTXnHP1V9OQ84DUNjRMj89kts68X3
M7mgYCuNRNM4qLEV6BKU66m5HpfpqnFux+z6QXCpGWqO8I61DAamZiC/geHt87qt
+zZ7ae/yBHr0dGK1SthYIQvdPg7SF2JKhE7YBHgojXCpPHzM/2yPFfxPHzlFntqd
iLlHwi7yGCQylkmzTK5OQGQ7SVd6+PjtYuD2DObBRcNRXDXtg08ekni2wGSHJYJJ
YkSau0aFkVk8FZKT8eNPm5JbiPkIJH4pMvMDF7Zvo8N12evzXfEQBPCOjS+rrFVv
QmJ9TJU2O3s4EKFosaU4iTsEC5LqVndMKRoy10/YTI1Gf8xtz+fxMXlafrRDRerX
w6deaqsLfkkHvC0q7LqFbk8h87LN4zQpyMKPD9m37LHWhO7sVj/cHFQW4QigYpP8
9mglFstVLinQBQaubDIKSjC6NCc3i19uV94GxPw1vRrpnKitbjRYjNJlKL6zmJQz
qcAnIC9H6a1mpY8is6hyK1111eZydAhI4j3s35Afg0pVKMAedHhbhcr3HTMDjcWR
G2oQqOMxzstR8vciaBzthhcSkZspY8AnUUJGHuhvYGhbP7FhEyTFDKixq5h+Tvcg
SRKPeNZqTPytAr1B0ZIjyffQSByxGOkF+sdy9R4NMly01a6ScSUbrRELtDGd8CrX
A/ks1aiYp+scA1eeJLi+OKW1+IAoL/NLbZrtray3F2aOgfUfKEAgPWZhAYFMQ5u8
g505VhmCNOVDd5dAtVO4m/3V3th9kuf5jbXrPfXnQ9J2PKXHsNVSrt/oVa/2AcXT
Ka4M7r0vl8V44cASzcBJilktd5KpoDwuTdD2rHzLmE9zmIBB+fHf/sRetMnIAAVA
m1N7DkJk5XWwr1aoCkY+hR2Nx7nNkJckfduRx5BSnMqKF7BOIaUeLQ5bVCB0Yfn4
LMyxW1lcFD2Bxeyco/TGk/DkGkWIQxgyJ+Ga+RSQoDQxs3v5+Hx/Nl1BFnn+wip9
sApTrCzQpkgDkbGo2z3NfSBcawoKhQrjnpkAbe/oo1JfiaQURicmPJakd3bA7qkx
dord70VxG7waw2v+113GoPykiKH0PgicERLbcNnRiXgnlNgRZj5/W6PI/xVWYpkK
fEv3TRh7IaIwJfE18DFWjfi+L8q+zdwkh+e3Uwljz3uMvkhD43AnIA93FgGsZ/61
SfeYfnkiynCTjq1FKPi58BOAZeMs32ercDedxeyLEm2iErN3LVuNAWDu4Fliaq6M
QGC/FKviAtHE1D7DERdDw70umCXLrisNK6dg+wKeKSPFc6iq5ZyGylPcl2mVi1he
Xc7D2jzZU0v/utGJr684NMOu8VXRJpwe2cwC8zHhZO6nDpHZQ47uBzarQf1GvuDs
U5o/+zVGJ7hJIPI0ruDTGNDYNiLsKIpmxuUt9BwlXF0E4EvTl3pPEDg1YIxU+YZ7
mA/Mlqj7py+AVRIc9+OD8nmxUnHiDU3gJRdNL+mnIfCZ607n0F//khJPPnIFqjNa
qXvJI3EPtLc92PuftBTTqWgc8foH3lbz0X8QhCpk80w8rsjpY/kufy05talDPJu0
RJ8GhyPK/gpQ9EasTegmygjkK58PturoJs40IUp90HCXDH5bXWfsWCCAhZVI7Baw
DlzPR5IMsf9lFWJndezPSwRsKevwGKu1jmYgTao7s8WW8XyufrnCwaFdQiz1rav+
0FEMpik2o0wUSX9M5U/5yXzG4VxI0iAyY1AsUiA3qnD1iObWJHSUL1KFvlqVHgz2
ji8txPZCcYjP7pjxVGdqfCx+1rSNRdNrJuopHADxlYoN2V1Qi8sdmWySwzgFwwAO
2JfgWhiCVo8YjNVjb3OXSsrbTj6a1VdRIkCEjkDq1zQ4ACkA38yswMA3CvZNS1DZ
ZcqCBC3qlsSgnd+reGirSq8FJGSpcciIPSW0tUtYawbfHvQyhhDsR7KYHTalH8TH
ahRqdWtCY7xfcXYTGft3oS2NQ6hC3bOSM3pohTrBDsH/OvRHMzg/hSdpvcW7GM2B
AqLjH/7BmzzotAQa0VFNhGjS4D7YeGRd7IyOWey3chK4mDf95K3idsrJH0bR0tHJ
WotLE2AWlNuHIhpjYzgzBjMXOLCg5/Y/3xq46zG4f61WW/Gci8iaqkqRMexnwJej
qSTBQo+3//Gs7aNWKhXcnh2LMLSSD3JEGHPdBooqS2mUEZYJSea9ZePLOMjqhfMm
FQwg29edWwYyYrD3neT+l05m2Y5YpdadmTi5DEzwLJBnuOmQ2/KZ8U2fFnkwOZJz
LV+P7WnqEbg5QAGa+gz2M+GiKnxfFMw5gn6oIApeqrv0E40PhHdJHEGUNxmSQKzS
5WhJa7jKg+/k3roEzD5SperAlqEK7+BlIIHYVv8ip0CNAiTV991ypCN6YNWTB9UB
g/ZHRakfu6HD/BdfP5+VfU7KF850tHDumsipIEIO0qRNJwadFjzkNINOIkY2nDPJ
36+SJ+ve+Nnr2hl9kTq4cUS9sAma1O+QlfNnY6eACaPJxbJIHyJiA2Zg9LRqDafO
9eDA565OF5PUs9wo9Ymjh7z5cpGMbbE/zd4O3wfk9AHjGJLG29kW1SX+R0/Vomre
yIEIa55414+7YUApOmjm7qf19UoyXkiH+2ZgV4Cce24uq656XE3h5JfmD3DQ8piD
Eu+fwv/nb2HFmuqbsVxEHRtnnMGyuWDiN1JDNvq5vpCC7QpEtuRFLe3PobCmuKuy
hdW5qNIEQOCQF4RCF9nPgjb4OoIonBht5EDQXfGqGC7zsdcrLtr4XvyP0PZGo+vT
z4PmOdFs3rcoHPporZOXFYuTMdyNeM6Zd9h5L5Ux1kmPoxfk5uEp+6feQbNbpqRc
UkhdLIY+UwWq3bpdmf6fcjHmzljT5kTs91Wfnw5kmSWuSKFsKsQ++dT1ghYlw5kM
/SrL0U8WRyeT7XIl00duHgxhPEmN1ql5NnytDR8toeBAQoa+G1GCyYuZQ8ukTrvc
Jx0oJyCeQ03MwUogAD002KJWj2k1YjvPlloPaX30H96z6+9HDcukLvDFVFtP4GrL
/9AXMi8aan68uUwUI/IawolDtHSTkwyF9AAuRJglKYzKIi1yctEgodfRsycwYb00
BBI/DyYwSJATZ0VFefrLzIrKshVmK9Td+PRfMOLutHheJQf9dKs7aZ0hSsOndKDu
siA3KNpkiDB2sy8MbdMn8lpbfSRwzAOeYyPca0TJIEWY5d1NvvwGdKmlkZ86o7JT
E6sN1sNoyMuC+QBgzn7bbGBQiithyiYw2Mb0H0ZhoFJ/fCZOkQQakBHsim4RzeVh
yWXj5gLhEFPqameAPWzyc1zqiU3gdrzxJV9BH794EN3oAKRaNVqKtKT9f4HnLiOV
pMWy3vUxfoArkdit+acBG5maoLzRP4HBs8y8/6h1uQxCnsEcKYM6/gqElXq1XAy1
0vGzWU8NUnzeYW15uO7zIzwLgoNKgU0H65FjN2RAUFvdCa74zEjxnHahODDZqjOw
dhWycaYc7JGO3rEA+uruif9i/3qeSY44CdxFPOGoSQVOk8aP30iNl92bfM63mqHj
JITDufG36joYxQB1ve6Q4jXJtRqyyrdIZezzT83yBAlul67r+rlqDA89JV41qimu
T2s8h5VkYKcvWg6IOuiJ72AClgjpjNWI9W+V0ByfgZ841VKTbavZbkub/W8M9QEL
fefmrWgDLA86HxGOev8ZzaEOn2iHaOxzATsaAoPhwii/Y/GhI41gC6UleGUKzva5
ZeA5aMcy6mlpA7t/w8Wom7B/NiprjrKtEnXAIdmDmB0zXO0qIoDCGEZ166s4nlql
GdU48SX9YghD2t79sKdadfhVZquJ6Db2YqxO/IHOEeX8UBsHNnNtYglu436U4itd
C3lYWb1JMBE5eIY5+ECyvkOj50uk4qO2qturOiETEtxiSz6/8gN4NMQGgkfoQo/5
JWYFF4CfXAHTXVZoWSWP3R94BoRONGsuWKVCqoeTAOsMeLMwE8iddW68IHDBa5QK
3zHFSsuS55ITNh1PCzWAYPb+Wo9FJW+pida5OjxtN94N2iIv/mWISnhXzpK1XoS5
T3wDwR79el5Z4Hy5ULPcJdw71vXVg4r6t4EpP4acKfD1dwkiZ7uRuX7datP0cerB
PZrSdHn/Ta5MF1C5raQlkEYPPlLuPQvLQZOcQW8HrowGxjUBy3SJBwSddTRX0eCR
b/oLkmWuS4yTpWpBq/9JNBZZz9Rcgsi0K6qDZYRITj6g472kIl4Khi4lQmMHawSm
tBFmdJH8jCMyvvYv2pYVEFlEF27xkQ6E+5039eFc2NR1WYbXuBcB1A8gLi0wp17U
J46K9ZCRbAn2MlJ3yK8Rnz8+bfzwZ2xqTKwc94uUWhR3u+EWKMCP2PE0114Pgaq3
1b3No9Tl0w+2awdbSl39kSi/udRWTgprhZYu9T5XSgGwv2woPbP5aHOFcBEjZ7NZ
e6rPwxn/775b1tKokPBlyyK6wMfwUTDBLpL55/2obFFtBAt5eHirXqaxahO1td6I
fvbOGB4e7COP0IpOGQ46Rgh77sEQfXC8/nu5j+raAkEzaDqvx6doXJei/6EOYALD
V88wQ/mY1ls94G3tJKcuvS8/ey2tZkdxuZw1U3KzZ3JI0iP3RhyNrKNcXy9STg3G
sw7C+iDMGJPL51N4T0LsAo5VE4G7wc80XtPIE4PNIVWIjKqaTCXIdh8l67lLDd1G
2D0/hs0lOgPWss5PtgFnvAF2J/XRzUQfNI5FFZoOaudUajW52BW7UOPoj+HgYLlG
PzPFYm19cwWsKkA27RfDKEin4chCTf+1btBAqiUwMuhkyUsNu3kFuvXDb5YDdnDc
1pFaeSWpBBifjoXnuF7Pta30qiKqARAajTDnpPCLOFSASikQR/3Sa/AtKmUXbFmV
i2RTGisXfyL+5RpDKLcHiO/ivIcQB2YFzP5vkYZOL7PHVfaPv+dAQ3wiGkbR9+UE
ecAR2R/KfLJJ/++HVMIWsD+VhohQpKx/KTY5cy2iYMekxVIdpxgavcUf5YxUQ5UF
X6KuyHXXjQTWl/tHDV1E891AYy83sZfkzteAe7fGDAd1sqxe0ZyYYjGB92cGshZ0
FNkMarkjizPIvYlulrqgd+bRVYCKzK0ZLpev2gL7zuLeI8Aq77VvHnzggRZ/sy3Q
nKaQ9f2wdnGk+mJa3deU1bGoMEh3rA4Pewn1Htb/pc6hZmjWbJcb+UY6U1GFYIkG
2YPyma3eIVUJUonERQkoPt2k9z9rzsvaTSEioFdVWkszK15WGyL3MXhKdl3e13JN
HBEq6VX7izVGWXGiVeMBYI8M9rZX0KiNftRxDKD7GAhS1nQsHbB9d0Q4W61A2VCW
9KfByC/vAQRS6Dky70IfsXQEx/lJXFyNi04J02W9ZxHA2mNSbhI5ik861plvtleX
hoTinthUiBDEwHY+tqKxLr6zkbhOMDHZZ08bRJeLlHR3rx/FxHrW0CufOHxuWQu3
RbfuqjWiFSe5It+J/pFMV9m5ERBPHhAVRPviE8/5h9HedrrIltgE8GAnF/jyJXJn
l15urMeHlPQiu1j/KOipSIVq2lsE2oh9wcubsxtksWP/4tNQdssYpA6SrpG2gZ5E
JkvTn0CKofP/cge9QQ/xpGuifPoQ4dJ6N9kOPO4EOb1KPgkYUAQH983GcjBrM9MV
enf83RdQeix/4bVa2XjCZmmi4yF0iax990HBe88EBQgQWIF5cm+XLhoPjT5XRcZI
DiXmDAB70sxkrg93cNk/AjEodti38GvvUOGFCYdtbCGGk9gtB/tynwZIZgGvaPiR
XJHYb6qiU1tSE2S9leD0sEy91JVow4RurQB5NI6wnHEMa0tb32uoZy++rCmqMkFQ
kgqzaUO6qHD+Oz5gabWinVCanAqvPgBW2XxX4WRZH6wLHujPtRu5Itr9tGM5qjmJ
/n6jMapMqwgAQpDOv1q0JTMEeNLvS8cJJUdqKVyzvgWZ7AtvyO1YoK4c9ASLsYyI
wuB5StF2l41cheU3CLtccHIwtPACaegapPT+R+V9EDX1rXXtWbL/TeJETdSKRt+W
Wo6JIKAxN2waCllLbG2lNiI7sHnP+wH14Ug7B4POWXOgEBze1JhOBMyzizH1k97e
MriVSzT2QPa+6yX35ekqaklvdvvr0x3qEZjOmN7oNs8Mvbnt7Tc1beB4n1XjHUn7
wTLerk3k1squEIWLAjpTCt4Kyk7UOelL6Cb5azXi3/nzCFv0QHjOWY8EZfHTT1ck
k4KV1GDU16gCq6mrs0n2UDcWc7kxdLigNPToIs5hKpS7v0pvn3Oncou+Evz/8+qC
R5z/mGSnTZmlObJAdvwLanOt9DPZTxIKPXgLZLUaKN4bK+gsrCsdiBeN5YqpE7bZ
aWAxuMdyclRulC76wC9HwjVnp2KZrz4wYg1d2ws2OG/tECoPbDFBaINywdMSgQHp
Scyt4QA3CbDLCFf3v++94H34razdLCr3FjFsrr+QpiILTxzh2LAJv+4FRl7pdo64
egzslA/0nip8APL9rmibvoN8s2bzs9A5UxyugcnevFxn5mNjPGSGL9sHu9u24sOG
VM++RjD25/fsfC0nrnhsd/P+EzZa8jJ7tjvXxWfgjkFDHbnIt35Fj0MvWJuQM9ZX
wM6g1xzSkPG5LbD+Q/aO9tcUGayzNsjihR1/KX6EotFqVWK6S+ShJhmRamgrIAcz
h3zvvY0+VoabGcycqYnl9IWz1GRDL+qknr9lIe0BgR5vLgTt2lj4e0bljKF4AyHv
Jwdg0D08rK0eGaDvlUYNGEyaLgWfS6qc3WubrXX8UsyAIGRThedDT0Ctwl0LxxtY
gHuDGQVuHfAj151JqUOXwbWE1yN8g4I8qviJ80U/6rGOqXYjYB3gDdcCzq8Rag4x
fvaLDOgQMgAkr8HHEcS2DE5XwPdiH6J7psAW6Lbr/c04IGvUdue+8R/2vtkCQ+oL
upaySfTI0OWPpHk6/xG8WUapZrbufzJUFfaKZkCmivpexwGBFDzGFJajtLCIBH0N
XtK2wiOm6ZgAlacRh32IKPa997eyRXKPymDY+vhp25MJSmXnhQ7ZTTBXaiHDijFb
9KQ7rhnMYCG2Omvuw3f0VXfz4RuwoBV4dfkKVMKlbDPFdzFYuHSy0s0ABxsgI0DT
i4VvA/mEeOzM+3FH+XKDFb/7Zv5leehS0f8cFRV3Yg0VkkrNESklU9T83N7HFPhD
oqpKdcsPhB6YIW4y55x7URPpAZYHFJWHDDxdUYFH9FC1HF560W6AK9QbKTbpw06z
fe0krMtcOb85/ONAyGc4/Wesv1+4aZUXGYaOsQ/VIElP50N4tK1nNypkUzcFbaWr
BliFGsPR5arb+LNIh5Qr/3GsM3Ckcf9NPrLgCsIOP5PEFzGF+79VtpauHhpVR1Wq
k4rrKSlDtWYNLCguK56JFo9isbnHHak3G5vSyfz7rcuYoxZ1/Lt3CtOcDuCGk/B4
nGqUOFE4PAoZMNUFfoPCtuWAz3lkGUTg7hMnYNHNO9SyX8kNSNL8WeTDcgsluGqt
mSKblVbfqEgleOvVH7N/BVv/yfvkvOdBc/UydGOHd1Th9079VpqIPW27fWJpizUN
xfsvbpKZzB1XVVFh069DTAf8X4Wpy4Xy7tYb0AXmwrZsbRPAOPzEyK3gaIiA4mnW
eOs53cJJWqGzqQWlTtZZ5Z4oKZ8+M3wru6ChdbvRDjkuThJ9KLo8FWBZM62bn1B2
W07cLf0s0A/IY3cRw4kGPGw/+mD+h701lrhmztXqCHsTAY1wBQaw+QDtpywoBJOj
GiwZlAmeC2WAZZCfHpE8I6gxdDFyDIfVLX42gG8Y3A+0Ze5Sh6qNJQxhpV8h8of+
SOf+4dMOSp979ZEN6a6hV0CgWjOU0ipSqn3W1dr7J/QaJHa7HMjKCqD6kZ6aQUgT
BC3LwS3wRq4LOo33cQmotwAwedHgmZoPtzk06/1TYHd6I0ZgqU7pmapSnla9S4yt
JrU5HlV0xyWNweheMgN+hzeZpuzuLckpv7LcJPQgNcwVKk/s8S//yDVdY4BEjC1K
rKB1f/EygrTt/3Vm6DyD9PIi0fQWmz5jYWb/G81KgmnY03f0t1vcMyGHBmVxnP3G
CZJcNa2LEnPTCCJ66NOTvsb5DMhCXlgireESdB89Isa4q1CSiKy06EMuEQvhU6nJ
55mrH2M/OMAA9bl/CwGiFovAHfTJQFHzQK/sBI4ZwLFjRg1BFR3nt3JNEdiA2npN
hBGjal17m0MWVDQh4qvpmaytK7fgA/M1s1FgmxHPwxe9OWI7Klv/lc2NqQYaC29u
0ycedRmgLXNtpD5Bsx1vbdLPDloPe4ZBNJuC8TqPU0QVErqrbXk6Nxe+bXxmPd/u
CZRHVKVZ0n+/XgTrOucjPmnmk17BNLQNKtH7T8/yb4jPkS6WrHKFSwWKrAavQp/b
UTgsb3HGHiahjE1na+MlCkg/aKj4/ZcR9s6EQoi+pi5Jp24wIY6Vj7JJ0TIRUe40
a2hKQYBoB6SMd8H6KOxQwRyGWV/L/kJhKQIASGbjY7ub88cMVUgQazkudEe/2woB
sGy1TXbWmp/XdP/SgJtXWjJPkRWIfGAFVv40KdgvsGfbZQldaAmapE3T8DuCJUNa
0wcLtvqhNwhwucD1wMpRM2cx9vG8UkFsBWrnF/3lggeFDZUu7SJmOlfOaaUiy/B9
HpiRHRMAxXnipEtfme5YPRuM1THibckZz/olP/VmQbxh+6UcuqcGB7ne81J0frRq
9BvOG4MmCjKD6ZAwrRyNFQ6t51mTzywES1V4Uj+jlNT3n4P4LMF5hoYQPgkNLKmO
HUKvut+4WSJG2kPVXdIH8VlY9Sc1fqmzvNQnxqh5a32zW5lsw0vH+KsxaY6W6SkJ
5+mK7ils33XnZasRQ6MrnLCN14HSfV8J4u3KkRMMSY0IAW9BK05gDbkmqRsWaicb
Swmpgjo53AOJJedMIdUvMOvWkhcfh2AVYA07FrwqZ+tWe1mnHgNXkk6VsHPGfowE
pZCzuNY0r0JSW3bkNkmy+F45R8/5RwWHk+JNw5BJkjH4wz1q46/rliXjMVLi8Yw+
5Ij9GzADpUMm8iGdBq1FUQ4Ni0hvGV75ivWhctXnuE6uOwtLl2ZDbdTtrlv6shyt
1xwSmCmSFKrDjz9k6EmqsXBPoOHBnEmda82BL9JoEBx90rE+YXh7gqFFZr5e2wcu
q1vs0WOFcO1OBHFuXZWoj3FwM/pMOvlneOkJ9pbuSJ2SuCKa24rYP8iPyFPsxDKl
oLpeY/pWH7Pb3A1rh9cDupa8BdW3+abil5KNSzm3DTTKuUKGbGla9NDy52QOgfum
6rQcGb8+MCxQLaGSm3Q4Di7RLTAwlpF21DyJ/pIoxXbc9w8Mm2r92KKCtSJQneha
jGX2flVVAO55SsGwPZB2Y+M6SLMf84HWftZ2DpdAyo5moMAAv8H2PEFprqJAdmp1
FyfV/MpZ+maenI8khuaa7bkhT76yBStI4FuyIHJccFyosQw9tYeCw6dga9WPpSOT
jCBKqt7MD881BcF/s7zdJNmHTxj0f3IYN93DQUjJ5l7GXUA24hBOauIwv8Dzf5uG
gJh5abQx9NZNO6OdUgjfLHpbb0IDnKkwwzalZokwCszoaJ3QmBIQvKUkYkp74oGX
kNll1fGTqaDFa9tfaR23qB/Lp+ecH1gw64w/wey+KfOa2UrSISvLFGT5452oydJN
HB/wOpfI0h/HfL5xJjcUje4tud++SPo6EHkt6jKb70qDMOPECFkQYUwHhoS+KNJ+
5dtwk9EfteXC7nRFUPyWpLmtmtFHNb843ScMunaLTl4VAv01u1O8FbkW28UGO9lc
xvOEuzHWR9DTI7e/eMJuecAtEmQLLivTdNX/NUtaHX0Nx86oUla1b8CwtXxtlRdO
ATtu56FRviCjEf3PLRNw+MXK+3LUDtwdA4nkxMwyIJzEeaRysnkPykSIs1V9TlNA
0rsp1NX6AlTdKwkDT146U7jlyG+NjlxNMJFXRcRQu92v7qU5VVpbrwC/Rx+egavL
UFdnjVl1nsabYpUT1F8JqvtJOapkwa0mcn3ei/VK0MjCuddinLufIjksmKQ7FY3Q
E4jxLgZJ+IUK3W8D8UYp4Cl58b3XWM+0vo3iRfWPwcNOacTj6LBOJFBHqthp0fG5
5SD9qXVbbIL8t3qJVvmZ2PCJ+xcvYhLPM8jNfftwiQOHCI3Arfi6H5O10hA1esJQ
3VkkKRrVYEYxEWKAV6y600qTMJ17mB68floKvJywvp8TSxajPb+uGkmEw2JmVT28
GCwbc2zihgK+qO6zlreivU+31uWbcyyCAWN/ibW5XXxMtvPi8pJRKpggOUWrGuLG
8ngRV30q6GPPEc5FdPrFuC8R/8DGXnAzdicn2mpQ0kj7q8RkI8eqEHELNZ1UT1Er
6XxNv/7veYnnoA+FFUoPBjQY7X0r8vphGZNjEOxgenTycygPIbZ8QdHcVu3SQbLZ
5In8m9ClyMR3tjnU6GZZ29g9KjKrtzGwdUiq+loAJtWgvr5Mv1JgpYtwtBgzM0s2
NJ+hxHGUaXNWkX77fSyPBfsT6m2H2WL9EmVLc+X1VvBhq0CzNs6+zUNVsa32svS2
11+LBGSP7hI2R7bF8ulxxkWvpYiPls0fV0Q4yq+5BFY+/HmCyDC9/WwfnSQOFxWV
qshaueaDQTLVCXHHnV0O5elykZ+/YqNRRU0kxkI/SjgSwC589/sEjmIie8vZz9iS
oRZ8yv0I/CZATdKQkC7Ux8vxHhBThyiu4XuEw9MHtUT3ve11YRtqrf+QkmyrBgME
CB7qgppE/NR5rOl1ewcR1pJ6ilWuZSd34+tJTrokVgDM/WsZ07o5apBuS04TfAYR
InhSMBWeycpaQEoYaEdqWwM85Cl3KM+DwCS/UKGpPuBI2wm6WLkM5+cPAFXADZSB
U2pTb1y63UASVhmw7y/b1BH92mPx0jZ7UIgOwb52245S0HzoJQ6lg3577PMTrLO9
vVorjosb9socvgzEeXYJpvIeY3X0JDYJpvUCPSswEULoJe4GHtm+yAi6buMt80ir
TkygdhnKklRx1x4I2ESn/KGnSFAbre0AjOsyUPKTaeBcCEBsyAsAczh8MqknEcHd
446Va+MWF7CYNO+4uzcwspYVhOMVSO8A9wjtI2a7O2ATdoouvcEB/BaFfIz5T5vi
ThQJXcAzs523xpX+3QOq3zLfgdW7yKyecL406XiAQKnjYulLPgJuTCJY2AtLFMIj
tR05QsaKqIce7p87DC84u3yfGRnuaEFdspy5lSXbVY9r/RnIct7BDWVNSF2FymTv
7rMvwWkc3al+3Swc2tGP0QWh4YP/cd42cr52CPcKpwBuiFm8V/aLWkbLTGshS9/o
otY+hLg5Wd7tgovDB9m3YDFCa5BBGEbJgc/jajUG9r9AuisuquCE/gszCWjnFCyI
duyKP+NEwRAqSGmm/CNUpYUhZc5QJN0j1tRwgjpqIIXxGanvBhDhOrbyEIWKkKr8
/mljErRJHAsfk9VNzCuZPxAWnSRYemSsc5ssxci4ig8YM+N7mkqQ88ozSQggtlMe
TaC+obgYhT/yXaTOdyvsRAu2cubbeKh6sYz9YmXNXE1Yt+g/mdf9MU3MSYQRghqw
F6cDxL9WOqw4fT0+m7yjWD+zHnP79yJMy0hGB49bqYkxN6lQzBgxO/q2+lrD5pdS
UVVbRV9cnuO3yUDtSNV8ow09b6sh8lFaj4+oV0xdnvkdr2mXptn7mecEFLvKB/G0
dfltp28aCB6Pm3kro2Bk5U9vqCYNKbRghlIcoqnkfHk3akUCIvpqQX7FADCQeK8W
dXuapK0JcqstdOY74Y2sDO98LOPH5gprPKClWZMIhDp8wHnIDopxX8oLDPQsM5V5
xP3ahCtFD6QOAJ0nvV2F8CHVF/r3f6aIAzEYJdfgVxpBuqFb9Y4QBsUAU4mUVket
yLKjAMlUFl83B91Tgh3rzKpuCU6v8KgYvSaXoAVbuyRvbXsrlkVT+i0010WW5HPu
v4hGv1XAEPFORiFyjBOgMvcFHRmYWXW/2Q+RbZk2icEiPOc/zjZsjUEJeN4osSmw
zzjaFYES53LWoiT9p9NkvCuJGjqmdziG5R3Ivcqy4EaOX501e8T+exG/dkb+ve9D
TdZgOxu/TRSS8g5Gnk/rVfutYpxhKsoF185zw2F8xX8niukD8K0makD35vTagqYB
VTPLnTaXICabqB16by0k1KDW1+7s3ikTM3gr3Vr60AzNmSRCts2hBiwKD9Z/Y4Mv
/OoiPWt+S04jtQsXeBuVAhEeO6Z5nRgXw4nu/+kxl+Jq0Lyvx8YrXSImMQuV1La3
qnSBJCD1bHX/95QPi8cvnQvkayF9NUSV2+jhEATWEdFZX9K46IHlN5Qnwq+bCVY/
JZJL8bxVyV7lZw6xNmqeGuaSJ4NGjXHAjMEKtTxDrtI4ArdukxEvcc1sIE7IJWLl
JMy4V4sJk3NjDQjd+8Gnfs5u39mypjpTFY5i5ZTOedEU5nhRngbgj3v5Tcyn0PNk
+Bj5Y2c0n4OF9euW9uYr+oJG34sA7jlY9aBNjUDjaUks4LsMOHxnIZMDH6rDdAEu
UfhAoL/jhT8alKozvh4Ujf6fWQgfQ2muMWv3u2sjfBe5f5DyqvJei7QUp11IHvhC
lTLjymKmyEAM4leqL1c48TQ0HBpZ3hNT4GXWVtH/z8ZqbmZ9g0svNKggiCrDWs4I
+CvbzFmg9dmFfYaOIARkFnIFWSHkc5GljP2hade8AoKtw/6cF+S/3boKddEG2xnZ
mvjJqoAQFuTngzEcMbDsWIkYjN7W/E59OCgXsvG418hxkEGkJT90+G/pncuv+H4z
j1eb5HeuatB+0ff4cL2oQbt09AfsuQTUdictw7MlYJuaoR+yg/dngaXQShQ8zXf7
eBURdP9Af1NNDruZgxI15UhTXU9/QDILrlskYQ9++/zJ+DHomDh8nSFXneWoJOQz
tJyfJja2X+Afw1CvtguiVt08M31ZagpbnVmCBwO3NglYiNckTIilKnWTrD1SFPMJ
tH2EtKXCX6zeJWsZpwVz4iRNk4K4u2GGMND+yCjog8P5jMi8cgBJ/8bKkmD9t6z6
rTCKzZOLkpigytPAPHzxmT1oZIGMWfnM8Wogvw4qY+5YoOFOMzDGi+jtxTq8laNI
yNx/5OTxvQviAg4VKtXb03S5cOjTHCqBZ9kJdVYlSImKDQ1ZNu5DvlEZ3rYuQ7S7
1z5E5ZRjJ2S0roZhhzUnssXa5qBtBIqbvUbvJIwFWbJMPkLkB/IgCD8TXOD9ft5A
sRWRSy2xSgrXE1Nzeoti9aYidnU9qXyxRgQkzDc28qdeuw7+Qc1qjKfyus1ypIy/
yObl8vWddbkSrlRGIHo34Hsz1iY2R32rzj2Ny/uiBJ0ApOXsGoH68XPYt4rWPrRg
9pWDsbZhvZ44ppC2ONdk7Omn2frDypldTAvWYf8iK/cyZoTJJxjLZJGInvYi3nQQ
uOxz2SY0ZOoxm3oXAgBN4NRR9M47AiseySBZ4AaM9LpDBZhpyI4KDay8NW4CPadC
MHDEybNUcXIiW6ILNrm55FriCVcpaX/UWjMupnTu7Ykk91+zWLGJ2fyhUEsjeDtD
IwysXgQ+Hhw27WJffu89BIB2P5PTvfhXT3J3w8RjXMef2GR89q+RzEH57K1Lw/8w
iHy9czm5wmuXXNm1gJ9XgiLUt6yg6mH7FhkLt5g1egUOiIyKG2LNAOIgd67qlPDX
fj7CYA8DAtbvj71h9hmjzuPrtbxA7aVFD4+28f+pXgzH/HVHgKXIyr5rZjtoMd8W
r2utgcrDGFyX1IF0mvwbil07iSRMkaIA83Od3CsTtjD/4088CO6egfE2SeCMGckv
FHahY7scwJAvEdj4uSfSHphj08GlWEECInBvmolZQzwVlQ/h2GeewiiHcGAQw0zj
XaMbhSli5v1TaW9AiF9Q7d59/cuRQWPxxP8t3Z86WUPyG6FuavddgZp3Z3o4jC28
rHYoebC33d1pMC4cQf3j4oKMhunYOKbPI1LvWNMvA6ovE7ov0ih+fr7MJBcxbvg/
dwEuyuiJwEx11bYB8qr0eegEQEW66TtG650vbQLzhHOQh1c5JkqqrM/FCxr4zJcs
6Y4ZilbDi9ldqy08KIVbu5wdSFlSDGUks3R3iEJqH8EHxUvXKDIB/XxEFdU4ysG/
zRVHBJtc5oWxHIxSCmBs6NsmHDC4wHSqXrZbHxDauyupkuGZlm9/wnw2y/FFr4MZ
ZWeSB2ElLv4ulnscdpy5yqhHxF/d7uA50yyI3Z56OEmqkVnecdZ7gT/7egmw/Ahx
g8fEH6ZlzKQaZ5cYnXykXrh7DxVczo9JeJ5g49Wu0YcUF5yLO0NTPZkAEqO5oKBq
/skSr/k5KEKATkxkhXO/5iYkAr/Vcz7daM8jGKuNu2FaZ8WA+rdgIM0TZGHwD5S5
5fma8i8xXRv/P5z2dFxaIV+DazTIx5JtSDwnIGoCmTL7sVeWsVdSJ6uHQXlCx9tT
YuF8BegMDX9kcM2Rt3rOf1bjRsXwGNtsrf6TbkCghDrltpxfoIyUJ/FTwhzPKe+V
dmATkjpLGclmnn4QEVjqYTz+aXgmx76J8eGu9T3i5O0zEU06f9D+iEh1cR6uFzfc
A26qr5D7URbchi+glR6Ep5msWJkESWNb+3V1S7AkenATbusZNPgCwdaJD7z1D7+O
3vcvlYsgyl+V0HZ1a4murt85dQNNlw30c1avjdUqblvwygL6ft02dvQVzOwxr9Hz
0tQSa9hKMYtnxYhpw6OHb1a0lAcFVx2jeXSzx/eU46opgiCp9HPrI1+iOXoHwiqX
jUGDWBHPYC2/wUyVbtP3QosZIoG3/1S7ghmCKUzpPzd1BqDVY7ahDnnevEOtYPex
hU7BXZNUNjcHuBC4KFzkpvEG6bpabWmywYIx0ANgSEkYW84YCYMshArpLrZOnDK5
WIFUGHawRKIuoTDe1o0+4XKZfe+jvxDFwSiTL9MeBT/FD/2QkQNQvvQAzsXs1d4w
m8CS+AKqvZDaas8WyvEg/aQeO9qT5+vbfDA89Afv9y1sOEHjKTlbJYG9ujiVfFu+
veCKUT2/PfAeUULN18249HUr+3J4DNw3DuffvNXeEzgvshHWs/Fm7iuRljXH22+g
N2x1ejDy9ZMSq+5bECweB2dzOR7yy+k224QCodgrPpEIZWS0nBrMrRk8nFFkPXW4
y837HK+WAi5BdOJIVXApHDSaz4Hy0nioo6wSvXBxNYDNhKkEiTwHmq8vYPzcLt/c
5aaGxW38dnimr/4r7Kb9UmFtZYXAYlqNN7QXRaYqZz/7IVKbccl0QqeMB7GldQA4
pdxVU9xIJUHBGTJViRjmHVl6b+VQz1lp8rNew1kCg63gF87Z2FJ0ceUj8AfK+Gwf
QrqQFmvK5bF0C4ZqAVU2P7ExUQXjYNCL1FaqW2+NmBCxM0O4ak7DbfbII/beLt8v
lnDM2q7p4v8FHmiFZAUNX17n7l2tHbwaQOfsSZq/Dskkg9WEWmQgkLMkot4f1zl+
MlEajECjE0JKHPTOa4/n8MCK1SGVbGWsatOhsfhaNQtnUYoMIEUMB36yt0NL8vTc
R3OAPB/+9Ius++MZkDtB+eJZ3rlizwvg6NvIdi50HrPMGrtllgElCga/SRJ/LW1I
of1aMgsswU4z7bpgPf2pdQKLl0GKZvjfZEjDJKwFGDtUDD8pBoWdBmtNvQbaanSq
YCBikmaCWEdS9khKgpHxkxR379h/dtCBvH1k5m5eCP/IzSdMTXGgLDl3a/in6MPs
k1gGBl9voTTySntSnrX/BkjLsdEBd5t0vSM6feM/dXHM/sw0HgzbBCHfD+TFmmwa
RhebHxy4g38hZqO/1G7WvFYNT7Nv7n5jIRyZk5z9w1dIE1D/fZTp8b4EpYjRQTWM
EtsCkLw025XzkP0vZscREA4pZbFvM2UuGbZZIxaIHEKADYZ0GiNETPlVGXWZGcUf
ERUgqgJUHqxJmlo+s61Z6QnbSsIIByOyz7VB8DofW8OZPWJ45pabp0APR+kHE6UB
hgg2zZTfkkLoozxI17b9SAHFI8kEOfML8p3LPlqnbqi3wZRJz/rOksJFRA2BTS4b
qwEAo0bXahK400jlk9UHgWJjrIx+DfqdKsSuPQkbA7gxF3e7gSuc1HLjKq8eXLmr
vGOdhPdSMbMUB8k4w618/Gpjio75w6g7t2/J0hG8f/emNFfHlq+mPZFPFRmNmb17
xAGpzq4V1emObHsPUzraQn7i3SwnT4b2CClg6qJp0P0wPS2aLEnCTufamcsXWZ+c
PPSWKD9MaLRL1L22AipgXAh+Jcqs7ylpYTbDfopeXV94BR1p8cBkx22zeiBW6ldQ
af1c+vL/zK/iSNXqgiDsJB1qeQPUo3X69B/Tq0zGLFV+SqjzKMSErZ5i6X+dK9wi
MGRtCY7mIF+KxkoobVhyAz6BROdye6LmRVUB5bxM8E2v99rZGXbSGbOUscMbMie4
jCdj60KqLSa+7hTEpI7SL/MizumkQkaqXjjo28SUiLQJ4ZUcDeKCdBpOOjxh5Dme
tetw1PU4VVT4PQkTTixJbHTKied5r9K6Uyny0cymXiX3mYWFGY8m9qJmwnemsSZb
9kZlYTldUelWXZ8dDvMXAi1ZExJ1tt52lXcBRw8F+a5gEpYATJ6v1JQlrkKzMo9c
2plfXYt8XsTNTSMMA4755sfCr5kezmrKTnTpLys86MNrc6V0Bx4HLWp1IquOmrUv
9LEZn8gvEeilt/SrXbuTSoMUxkWiCEpDya9VG5oUvBZbuaqBVlP46DGshDT56Gjs
TKAywef1X4cxmtLcjf+8JNLFvK0rmzzR0Fj9ughXSsCNo5G5SEojZJZqnMcMm+CJ
ndTQgKR96hZ0dHshOK6YkqEVytkEXKsm8vMAUfzJE+l3BVeTqZ51TGR7BbZYxh8O
MuoS6o3+Zvi7BHER1qsCSBbjITnZ0VAjN71JdgX4dTusP7xVEKIc0cBV7Di9/9Nd
3jOOw42OZpVq4b7xDOaH4eBmJHZKFv5mZcMIQspa3/BhxEquEo33Kvd3WZqdSiJC
eHZ2TKk1hxQGibPY2Qf3PsaBIzC2sJHgF1ZiItYJhYvxs/0o7RN/v/1JVN+SuGJ5
SwVC7A/VJkOKM7LlrS+FA4SQwGr6kAg0treMyK7zNyajuMPsgNXEXF5u1szRs2Ci
MxM5ld/SXLRjNGx3qyRJjWYLWDu+zHPauqrdMoOIr2mcHjC6AcW/nU6+9A8TpTq/
KqNK+gwXSvabKdVeW39QP8ki+LRRsaly1WX0NIADKpFkve0LOFyx6NdRYKKiNEf4
eKWiXZBK43Nx8grVqoLiAxgPXOPcAhAu2VGX48JZMikNZI2lHIVu2fjuh2sOFg3P
5OgEEMtE28TAz2PvOb4KU8HWTm3eRuyeEOUwSwHO1Jrjz/ZRKTsQHwcOovZBfFOz
m3gSfRrSew9OMPrucIA5HbvrqG+UHhIBT1ZHAgIzTRwyT52KvSq0ZiU0yj2Dvvgc
aRbOIahtgYApeTyLVIIdxao0uEUOk6Wp2apGqUG16VIvARQ7hONiJqpU+uE3ObSv
rpkvefczl6zulEzjuCNEmZGREn22f6oNAiqaNwuG/qMeIwVNwMe7j7tjhe+LSzVX
jl2zWuQnd+KMrsneLzxKIP+Zp6UhPZu+1aFn1ICRuMlog58XzcAIDNfJQ7Uo3TTf
yjODZCVCrZR4/3LsdUTtoKDwcBKSzcwQP3R2ovdj5rjCsJtaIFqQAwnz8ynunmlG
fmW2nL+Z4aKf2mWLYo4pB2tO4aI+F1zZSehPOyZF/7kehfEK7ucg+4rnP2BD5y1E
rM2wfNKLEJMhE29DppESKEWx1P01vYShkEXYbN7cV4cWyjD3BIUgyXr1f29ueRw1
k2TfpiEj2c485B3qvKKLJ9uS8PqDn6NOB/IJ0uNSdoC91u4R4hiM954rIeSHKeRS
2IZZQEtRLN06RwxLPluyAwVed/AN9ZDSR/NoxF0D70xQrXc1kzBoET7+1a9NCYsn
UzqwGFvBK29tSsjN4GoXDPtlIb3AmGAQvBD5c8Bx+UFWEmUlCLniXwtk9lx1SHid
NKPyLsdr2Afc6zxiO5mC0Lgfv7sO81lY/PV6E469LixjLCsuC+q9CLz+KEZK5rk3
FCE6P/1jqyA9tEip21UBnRkoo9bWU2bsQg78IRtin0S9aZvkL4p6n9VzsnLPbkcJ
wA4naBzA9A2vGEHSlHaZJkErW+1VYY6Cp54VNZuVMDRk6QuTg+ZusxJ5mN5DHTE6
fFFx1qFNtnZC1cmlO8pamquG6YnjkoGwadS04BpRoxN+GGyxfATMfjfENSEIp4Nt
aisKhMMchx6LS+XKES9nyBwi/jQ1v4tLVb6TPTj/lGRbNKtPooKv58D6XyAQF/Gu
3FTND5RcGZCBN1oc+aDc5QA+7xH3imuL29l2MmGAzIngB31krSKnSHSTdUaAWdbs
W/mQTzS/KPOU8cy2P02D8OLV1f7HEj1mTnh51HSWDQTWxcn9MrR7T4BGSjuLAZKX
Sc6cbJPJ8irwyqADvh6M4b5ekuh8s7wAW+qMcCzmp4Ww7hgA0K1Wxr7aWP7QSIKA
uEJQ/ENLS/oQ3AxoeYchglnxx/AFTRJrIydkgHM7QYO/simUAiXCmzV/Q2mdk+lk
7E0fPdyKtJ59A0jP5MkujlmzoAufS8y5F3BxsBCY+vwG0eLZQBkHmR14eObHYjnE
Vw2tZz+uoBTUGz+LrP6UHa/CEu2PzQu3o8XiijPPIdnC9GmaBpbf2NaA9kxuXv0C
lC59Owqed3UPofBO1+HNMPZq1j7afHtn9R3RxT8VbvrdLnGqjExYlB98cBKgcCsb
tIOWnt3ALo6sZuK744Z8d52FfqfWUcQaQjubPsxvaLbaNov55kIIbvXjjQLg+FY+
Y0o/fAE4ViBiaJ+k5eYpHi0ljvyekTLBpAqVpybR0JWOgCV4ScrsR7dFmwHPEBtT
Bwuwn6Kxxe2IMNZvylxDDYBLQjmZ7UWrKqCMQOCOiE6AmEGYQTuv3+PbX6JuhdFZ
Wn5hVTnE4Rs7yCvgO2LTqHGMgv64ew40Ix2MIm98pmgKaSyjmHabAXJ54uO0nJPs
oOo5qR6V6bqGDUOsg9E/eOAz9BJbrki4s1tzgZknARzb4v88j15b7vsWBS/Ea596
xAMazMheUFZqsbubvP8KxqlO+ijMS4065+/Erk9O5NPyXjPOabW9WuK029QTaTu5
sWkddvUNYiLKCK37RxXMo31w7+I7FEqulNaj48npAlxS0LKlAQZyI8fvMXe1PkPf
9NeWR6eNbOPSSrPuLIQwcxvmReoLYCmjHRohV0TV0zlAvwy5PpVJQqZ2VaP03nPN
UUal/m4ESUPZbItnB/F12/4mUPRdUKVC/PTjfsQ0NRfiGKdzxQhH0Un9hPcR/3hQ
IKtk5+0Wm1jnCs7DcT0zzgOrP0l180CTphLeew4VGC6/XQIdNPVuIIjLyxZ0dXyd
mxmFar41gwQ9tMDxrHCdIE6UwcN5qtmPGJ1aa0l31kGK9scJnqZsW+sTYnsDcn+Y
AL3hyR82hi0+wvEGI7U+C0hfhT2FhMbqEvaFL0ANrL/z4vDsDYodzxnOAnScpreo
WfWFCpe1QSrhrNeFpsawo4wwW2Q+YccpEDsSFSMYiyyTa3fN87s6AYaIrvFiyMh+
TTUtXcEkB9NvltuXkp+hL1uw2j/sjIqA7CoqWzHWck5yfW806Heh06GiYig2eqKY
LH3vKamv5EyDFIi8abyFTZJjtvAt8P21jjbF6JkYO5Hd5q/iwG7GU13o4mmr4qwP
1KI6zRdovFZt3Um59qVKhB7Lzs8/CujhF1jKORDfaGRfuky79BnQsbGci/BfCjqh
TiQEF+vAsnqY4DA/fQy4fp1UgSo9DFnOAv7B42T3v9yiJUA1Z8aZngjLYalmbgwq
dbpMBOFZV6U4par6fUuPO3BuIAaQop5mtsp9qoFAO36KQXelCZpOvHrLvuonRhrU
mUNwEKM7vQ/fbfgFSTE2r+2C5xQZHLI+zn3OnVHSL/bYtlmQ6MKmyCAQebRD4qFn
uvKLDEswMXiFxZicmZ0TQTl5YQpenjl0gEzqgYXmkOflk69AHv73h3cASh7sNow1
mREdBbigPMDFOYu7B3izA09uQmhimqtzrQQ7p6ok2kDnN1uhw73Wb8Rt2gNCMFYu
nAkk6ILqTyISS6oPR3ZIf6gEGxgjCWnd40dXgbONq3eGF848tiYNP+GECCeVIkSq
moHjbVQV8TsNNpthUWiyE4gfVs6XW3/Jtw6VHHQFEVcfGsOCJHBSK365b8hVaC1n
37AkQBhAsOLHITB6pwAZPjfdfDwkLj5r3uWHUTxEjKniQpjnibnnnsWZcIfjg9mc
24d00nlCgRKMD5WATTjRRHuBl/qrEdEz9cBT8HSkm8zLWTfVYh6DHRjExRoG8d/h
QdwIa/AXcpwxtMDBrXHxO0ZldZmsfP9mMrHRNgneQ97Gq3JEZpiUfyHOIUUOM5+c
EQXlkEaiLJSReFTuqbGJp2N2VD4AJNV90eB6e2DxDCLirl+yP+C+Cum+gYwuWrFk
SfAgxUvZUABKB5QP9xS7zN/kdm631RouEKq/19bnUgCOErK/+/4Mq+ADofLQsAXh
WrN1R99DSi2SAwdemO2zz8r5F2BKWNbhZ40SySzJu43Ju512NmkGo0UBKtrocHPm
jceqGnX2Eh2lbtsq+q42DN7tovV9IazYCkxjfVxsYA8Ex/HKaoaOtDC39Yj37Ggx
QScroIklSMF/rq8q/EG9XUW4A+n7FPVikkMogOd2FdrsgI7BIwt8ZYfDNv2k5G5w
L5lNsAkXT1C1GTb4Vevc5xYx5A6R/8ZQ0j9XcCT6bJwBvtInHjE0Q/ew/fxMf8vf
yFn+aq1Z6oUuwQ1KxCtkSRIA0jpMCSYSVXIuw8Os/FVcCy9UPKzdilqcD3JT0mkN
f3sb7qslb3D9pZP/8E/jL9lHvvg+GB5jK/XUzNJCZB1bxjwOfYWrDfLj7eioleNi
XeOLgBrGcslnUXmT3o1FuiDGLVpb7Dfuhd670tp3p+GEWlkZ3xBM/7lUxFd0UnkB
J7uacXs8HlefUjm+UiZXdO9DzvBX20i3vXp0jfvTmFLGjarozP0m21NNFVCuZBxk
6Yu0hNca53OlqfpfO8JozXDCeEUwzDpUOMBbHBe4Y0up7HHiHlROJoK9t4MS4A6e
b5YPLczzn/fP/IHxtElPbQhKn0hASSWy6nuQCaQacJyVNPQE1E3zqHMfBmoaHGPT
d2HcXdWWdmvNYoJe1sZZJ8k/vHEJUOwMCw5pOR20D49s+VeJLUfnayPN+/nfw+jm
l130KdqbGJKiWNumdfKzyPWxCQNYPiGMkoa1mAwS4pLY/LtiTkOZlutrKXYPsRCH
g5Qx6KHnk/saLZYnBKlfJtGOpLZK3yMXW+/jBuO46zv1EyCxBZCtmC7QJOYgBs8A
TBiRmbw6ozD1R2H+1c3GDpbAxrqWfV/+UKU73ZXmoQwb9MD7iS4+CyqT2xT0/73t
VRtUNPE3Jb9uF1P+FXhunj7DMF+OnQ5VKccHkKjybHZwcnSejUqoKy6ZtotPt9L8
IZglQ7AZj6BBXao/srpGg2jjY9L5EaAWTx6VKgZhpl2SUIRza7ngLKVfaJ61fkpq
WLHY2xDG6E7EHX9QuqLmnTFmyXZs4gqak5FOrUndjVynytCDl5jwnDbrvvDgnLBv
G09Tdeu3J4IFDDsXgfWGNZBDfFHnqkgNIohFsEox7GnM5J7DI2DgpodMa/r6WLlD
Zz1qosxhF0BkHesIEm4jHCTxJu72Uz3UeWpbZlQzHnTpofi9l1eUKonnmc6ZSUjQ
divSvgPUak8/StEkQ1oHIwna2STEFYom9Qe304ODdkwtDLlUdhzZLWV3oz5iGrwI
So4WRObFDKmAVHyt1E+aKFA/SnFaVJCj/glzWiMHWsDw3vSN3oSiV6b6bRvb0Pz4
ZqKmCVQANQcjLX2G0TksnGe87TZ/H8pPAvGICYJ+AhnaRrz7bCuTWyyTRM17Y7wJ
EtbaTkvqWE/A0tBsf8kKSHoM4K+G2fSCbYm+ev14GByx8X60McfiSXa/zkJ/W6qg
FYfmMjIpYVrJ7r9vBTs+pS5yTNtDhzp1I3LtvXbz86fsI3xMzXZEKGqsRGlOiJjJ
loxH8Urbt0FzYDizyHBN6XLb9Hn0PXzppRTn6asZ95APr/Y371NwGZys9433OirI
TQ+GRGjOSy9OIB5fe6wOq0BUqtE4g8M870HqKQbN+UJtKKd8debx/MeqseWEsbLT
FQtZtJ7WxARoyT9tdwC3g7vq4bJmun0LY0zFlrZXzcvFNkp+swdxZaxR5Id7l+FK
/Quh4R/ipMKv/7Nxk9e4ienl87tAHVeFGMHs8/b07y+Foy6W+qtgqsVBPIz4mr+H
NGVOLzIAVzv8BngbB+iz34kZwZA54ETrc9uJPUCDKiuIsx/Js/nmZof7+SkRU5O0
nnaVM9A0FOP1aajqTSDewair52XrYTv0RwnoFoJj6I9onmcmDuoB1hkp+pyUSQoV
nMYdKT9VtNs8emM2e/atZ9t8XfDcYYamc93myJzi/olPAl27/1dqTft2y44RZC7y
R3POpmuHXHpWiWPFCjYsRfjZbu+Idl8RJfmcAnOYcCXR7A3TqCoek82TrNAyLnCz
npYNyvFAeUeHB8kvYhXj8ejvJbZeiUM6AsLDp6iYDCJI2K6cnjHGHfOhwafutE9d
gsVH11wMdefYyftAduJ2PaY8Gs12TbauRTJcIpJaK31our6tl90+IJYdGY/oRiBz
A4HF3KzWOY8tyVY/Kv39RgYfMvQ6XYBViOuYULmQH1CD1ROrSi+TBKVzKvgyi+hs
JxFrZeJKdgqCClq6zyHofrUuni3CeiCPa/QlqnwRmcfQENejt2RUT3jaYwTzt+zK
krRS4UIf1ck1qQd3ExU7aZ/tsWvuZG1DfHK+DfTIfFAkFTx1UvxzlT//KyeTv8Uo
sqxUHz/7DVmTTh3CUI8q0YAUXKV/XXt9tSnlJnSZZBxfXezhcQ3CM+zAJT6iOF3x
+qwpvYGUOw0T2YUdfCbPNbyA2ZamhQSZHElehn8rrm8LG1ZCmzBlDGOVACbUx+l1
oS7oalpZ8vUXho0dTpt+tzb6vZ7Ozgh5Mrhhlk2iXo32rJQ7P9ju9aKtFt7C5KTh
SDBPUEBB3id4k0f0txveGmMqY7UwfVi0FVEt23jy2LXM2FP+eiMGEmp9Nfl8bl/X
/1DzwbBJxnEQERqlaB2xEsmD03Z3zVKSis8S0QfYALjbAUgb0PVXv4Q+rSJ+cF+x
eV3T+cA55kWb3I+HsAH7WNwzC6UVE7RRGei7ZDi42D9Xsq1JuJrTe/NCo+XeFP+k
LsR61ucBE4bEAysKtDcH1tBnr/sjVuAwcNWwa3J1dMh4vXhG6vWdH8zf5nBSsCEi
lWD+wAVQ1fuwtwNTbDB8LtgfRfRnpZVkFqAMRoohaWNgwSRE/ayGHayJKUS7x8bE
tsSn2HefThq2uFJtT/hfWX0onedtPAN/bXcHbhiaWFqpc4tPiBl4iMbRozoJ267z
xKkTyBZ3hJ6rZoJaytxLuxurqx1b89m9egB1JiLKdGcjjyBcFiTkJNHO/MSWg+3E
VmRoq2RVpDF34o3SK5vyc8GNIlx1bL9fpSR3TtLDY6ofwsu1+T3MInrpnx/ZmHpP
iL9WxA7dbPuLk3MRlFpoa6u15iyirJ8zok9swceGZ/XLoOCAwRFoLKP4EQDFFI85
gi7aRaDT1D8yyNTbvzldm/LZ1IjorK3Zv2kaCI4g0y9HBu3J5DU0ddebfFIwpvdv
h1glCsuTf7n+LkWW2lh4I33NbjwAWfwekD/XVjuxj8k+LkqG6P4g9rUDS+jDnHEr
W+XhuZId7xChxpn+ywaRxGn/kLInAAeTa/4H+pbVXb55eCny8AEmJO0+e+KStJsk
43Ijzk5SCk/k1/lweNQgAWzADHSXE6vyztW1zORe/1xkjZ13jYnNvKcpXpsLin22
V+UnXNq99sR9qZ2Me5p8PoVXbuYqbgrmCXMtTZPaAm3fZ1Vv8h1fjBLzsZkXWLID
+zrHxImZsX6kqYz8IAljZlsm3cmYgt6RJcH1vAleFiXDP288HQYX7qbdQ4VmrrJs
YzlMuwxHyGlJ/l10ZsqyIyghek/wYG6fb7YxcElhnfvrXg5hc6ACCr4bqipH8wwS
I7lvqFOxxTsbx17VXZbuD3tkpEkFdA8yAWPVN1whsOypCfkZFAAESZnGmqZMfaNd
VO4eyacoQDbbVvZFS8MQ183yKnsFh4NbMhrHHiGyYaT1UJhC42iBUUzwcIJjKAfR
mIQJJR1/+T8iFy+LzzYcKS5eidiPvFWtyv2jKpzXHhlpSO/jwdC3ygvf2WkGvdf4
O5PzHnyPQp+fprptYpWRS0Un9b8XY3IQWR3AIgj3/GPSscT53jpkYNIEq3Y4EWSh
FTT9artSFQoGcnf7Y4GXPxAzC2/m0XhK+yruvVl85d0c3pcuyLsDIC8MoKeB+jAq
QP7qdZfcKsAKC7CyHK/y5SoYIu1VDF4VS25XUJZA+rppi6I4rPqZh2OhOZlM9HGY
YCOenF3Wz1q0H7UEa1qR/TP4dFNmXnfk7QPDSglHnCaNNM9/6UoC+uxscSdjBoIn
W/8qu9G7I7EK/K1fVl9a+7B2oLAmcDRGSFv+qBIkH7uk40NXpBU8v/LjYb5Fel3t
YWkcLh0B8jK2Y06BVAuFvsvM9FR1XiRXQA4DIxVf6uVSlDhh9akkWd2WDzLW/VfF
2PAv7+/a/oMQATZ9szt9MmTnpA2+kCVjHfS/Ni1B5kmameMbTtwMeG/zuN01uGl+
B4696wsWYK/ps9d1wOGThRct5109tRjQbY/ssdbGyeqRJA0gtWXU4BZQrcIFCoBb
VLX6YwaQyhbdjE5RWnQKbRjY6DD+rrXlAutyS6TBxWuFq/vFFf7DXaCuaMH/i94p
/G5f66Y38FbVA1M39eyvQTqtbTZRdrS0nVXMRLccgEVzdrWu8p6xLyOmeKhkc9z5
z4rz0YuWbZKFOxLjzTgpR9cP3T25KpeL8hz6vU2D80mM/VzvwAiYQ2XFVKF8shmI
Q5acxWBysV6AF66CBNozD38/x7egm00bNRrtuQpP2Ska6d2Ycbjp7D1P5BpjUCsH
i+48wndIkNPHf8L/pTSQPplX2ASuZ8rFx8ZbwunYs/d8Wl8zR2f0rkleHT3Y2h1w
X5GQSTflJXSGNfWRSByiv7Tnam8Ixev/ZfpxTz1daraPUiMLs5b867ZWyrMrG8sq
O8SLn5BaY8hUnbIY3l+g0WOWtxaL9wIlCrcTwaZe13e6F6rRGViVcLdq8TLDbdy9
zcEO/rvL4LEaBNTzoZkgtytDMetvWwC5+qm4Xg4kix8mI5/cStOuKf1ksiCyUDsS
i2ucIYStydHizMpuiJdTP7to9XPNde/+B+tJM0vcq6n17LWIz+uSqZ5XOLLHVu7I
rRE5Ve4HsY4MRP6EiQoG4P3GAhRJXf8WaOUGBupuNYDVp3SHpK33dWyDcpKJoW92
kAS74PRXuLwTWEPZ4rEAYHjY2vqIcXUe3GJleIQHKPIrAmFFMYwgumnBOQ4Tozll
3HLB+YY7Z99draWTFpJRp4IZu+cV6B/boWHiPQTPwHPetgTFKgNiQWTwacUF9+kO
AdOFQg36GvcTArNi3ZXqx9BdqhtarB5nEKcWEgyCYOcmWJvLbLbvnNUPFeDVkqwK
u3uwKHsufym9hS1u5oxisR2QDgeQiPNlbxEoLSZwlr7+oFjlGuqVomfZ+Aa9G+2s
6oJoT+ZP8MH21SydaFLhRHg2EmKz+k2mkZsI+WZtXdvGtw4hjz3ZqMBDHqr+jSAH
0GIhFd/51f4mMBgK0569qZrDG0sSLENK5Zz2AtBZXzqsiZhjU4LLkapU/Wm87WFH
Ej6d24t4C6Rah9FqUIu5EtLK847eNmknsTEzp0nan1Dx/XT4x+BP9s479rtChjFw
dQ0U4+TaTLMDgeF5VT14tqcSQmstIX8ipE9SCTskqSePJTM4oaTh8msouj0Oe3Y+
EKJJLEaDEDiGQYEVz0xnpZu7NjBFLv3qP75PdpYmOvKDc13bSH0NAAFe5uICKUj9
sEqD3CYfMNvmitP2Abv8tAw4rkeZ9JdPclJvStLyUOHgs1XTlP6Ml8edg8Sg0JbG
rJKX0jFeHDBmMvZmoPsg4QK8q3Ui67GQDQ1rF+82D4/6HNne53kHqMQS5bW2ZT+9
V8XXAchwR+VJ9JtSbJwug3JK2lvaQzKF8qc03uDYHtQbtVyk1109UGXETlbuMtwP
vWTFBPA+4NcDhwoQ4JCdOd5Y0QrwASfy3I/ptTovBkQ545sBgkpL4XghILZDGAcZ
6xwI2SXXaZ61gIJtncgyFwqCUA61EfqpEej8TtWvHF/YhtHD6Vb8xNNbM4h+w0SW
IYQ6/Pd+82r3hf42gmKFCJ/93NzcJxnUTzoQIiHZcfvCP0a7XrZ8MayyPQ2iu8Ts
6TngYzVBv73sdcFfpjcz3FUKjur20wS7dzBaHJhmIppqfRJbQ1wJMKXm53p+wuIH
fLrkYfkZ0HJnRANRcPmCvYtdyhzCG2vd3RVm/HZIxR1RsSp3TF6CoJtq3KJnXGru
4BIgeYbxFBqKjh2Il08BQDoawM4Hh3DwMY8hd9DhI3bhs6dvWxvc62JK2/hY3F7G
izE240SZj4u0udjjDF3xhPOqvNE9ItSf12autXtXd1U2b8BAFdSjDxSbXGXYuC2U
4vSHtXw92QrghmKGwoV2R7K73CWZV+Q+L6qiOMDveXvb4IF4ILDmXteZGcFtmayw
SOejD0qfI7K+gEUohwAIV9usKV2hJabeovuc4SEosZTd04Dzd6pGequlpM5wRmSW
XCk5BtlUhV7vUoFmTQDcuq15M42tUC8oguFAELVGANfkzvqasFus/9MF9K8oqTjZ
4UV0HL6KmKcHE7xE6sQHHup5LfbrXlXjlkxLDREGLPrRQyZfX69HdhBurZvkoyWB
mtTdXmawCFmxx6CoT5L0NCTGRMorpUSAnzGGU24HcuWjZffWa31iKbivM3afjDvk
50+hpLY44HsBW4mEnRbYp2tyNM71WzI5OXiJwl1mHwhJ/l0THJazjhyFEmnPUyHn
8m+o/tM+6cs/ywjEQf/clv53cKVHHz8MEhVDIBQmRyOnXrSR+lwjJykNx+Gb4M1z
vHodv1SO2PTbL9ActknHTPUQh4VxFF972x/RjipB4luxMi+NOo635F5lgIC665FZ
oJNAQGtMBq2WJEiL6Xz4OMOhCTVo2AQoCWPbkrSmmtnVwAOFBmRZ/R7Jef/uL5Sq
5+mOkEJ+bkz5UsAESP2jP9ATN7uhvZAKQSyeV7/NqHFt3RreTkfXqe3QpWOt+IOz
Ny08w9K+/liRTeA93vHccSBs9Gfxj3XUCtCZxrJgYnv0Tex+Wi185XtIZug6YAQs
eTnE9ny0lfesPAwzC5TOId8IXvCyQx3uYLp6PLY3B+OWFTcnnox0DlRObFF4Pnq7
gDR7w0dLBAAcmOXB5HFf1KZ5tph2+PqC6Umyiq5p+/KFfbuYNKep9D2qNIbF3FvC
7DcqRNYPpz5gNgl80T382f6oOHhw1Vv+Z28ti3C/7jX5RcbWrYsQ1TQalPYtE78K
vzspyazcm6Ynka8rzCC4h9BP0mSzubtL8VXESwvegylfHQ4EeF3R9ys0tN74dY3H
kMlrorzdb3iU8nkGwHvjMBFJP11CcimAZZ3Nl+lO3ZiCYNpeVybyrgr8s6rVJLXb
7LMCwkI5ss23hIcQnhyNp7zUyse4HYjlYufCkZDSe3MiIMZpSM5cSBnK4nOmd2AD
O7SWsLODIq4MeoQPWlDVyNjRrjN8HkFKv14eZJbXzpMHEi9FWVAmqopzF9PBweQF
M3p6w5xJOvChVIz3tAdSDR5DqT2KyOTniK44sJQm1Da6oi3z2msXsiPc6JSpqHT5
yCGaeGkenUKJ5GjCLgN6UmqHu7HOpHaGriGJ1l1k4QMfXUTeomedXTIIwHn39+AG
50vk8+IV8CQT2PuxqZAc7Ts8bYICdRzZnWRNbdfldmr/j+doEtb5x3gNAS2RwJYN
yvSbetseqSLa1wZauPrrKDiK3xeyG6959klmkhMzbI6LzMaXR68QJSfQvHQ7znNs
RJ2hqDpEq/dhc6dhTMnBJd0SPEYFO4odpO7r5Vz672OzFxHR4lef4+PQj/RNdM16
rXJxlIfLd9CNyw2jXMzjgUSY914+PZOjqaMwPIGwcAzJbbAYvJQ6tq+UOzUP0etF
LZFSyS3ujN0ikYZjlkKa8JUoHmZkoVeO9Zj5eVMgFWE2i+fjfw5Q93E2/R59OE5J
6Mr/l5VkKDzI2DQ0KTD8tjaKDCR4c03FBPdg12vG0Rzq0eZXRmN9rHRZcRe6Zypt
YO/KW5V9Kty3gUfY5hpU1oADQFsgGeKiXmVCXh+uFqsMcvXfdw5LOqtAJ0Y1vto9
a/Ev09QwoKXHC0S3w9hWva0+rSQ1SyTYzb3wKYlHVKrxfoc6Xpn+tNnBWxUKrrng
sSPJOx9LSdNOqm1wU7SQ3oKC/JJ/wQ0hMIY5fN4m+oKeXc4lPDy7qvsl/nJmNkB/
aDHn334ZskfMqBUz5evPfT1PvplRfKmaBqLq0KZ2rbm53Eb6ZoGJoV51D95QrNiP
fGB0AtRpoMX7OlyB8t29AAzZdL0IdhB0r/TEZqVoBK2COG0/qdullycEK8evD51o
gOi95pMVIOrOCHSTh6sEH0ARPxWIRkryzJBEbhVI4SG0ySrFCBo1oxYk4BfIW666
x66r9LLV8A1uJ9oYzzPSuVeXamwDPtVXL7OZma3WfJgEodwF22iLn4LESAJx3n3a
adyTWkKGF0i1At7+Nt82HI89RIf0w0rn2eefhkNr5LrE6P7AP201IcIS2s0Aa4Zj
wLxVC0Nv81wCaAvCbPHeZQ6JjHzj6hxL7ReYclnu4yUtFCGSqLAeD6DrDXB/Ra3Z
XiXWqS9Kja7o7DMZB4i5uyDRjeylkIsrmmiBVcaXLYHIhF39O2bpIGrYOU+J2vhp
A/r/au+xdRqfr4bULxg8UNZNlX2TZMBHkSjsuGcvAvil4ZydQqhIhe2JFLMPo7iT
umLRcbWcW3YSfCSvrFT5lyjJUVBplS43PDrPMen4tBJMyCSM5YB9Cu9V5VJyvXG7
+XawTuafr7v6bVe0X0E0iGiASwsJ9oRYHFOMK9HpTpz7yUpePf8Rht6SLd69NyzX
g7qAsrtjch+yOiqu9VL4l24qKwYx4nlJRrdiMQmldJ1D+ySML51xizr69AFQyD9z
5TfeA2k+Mz7adWoBnuqOknWdMKFtV4fD05CDUYuIltVl45S2WqOhuucoRAv+2i5v
Ci28zZSAZwJT9hJzwCidyL+GWvDgXdrMWwKTamNjFKmyuSBF+5C3QeDaAj5fUwxD
55Khbpus7fjW7kkAftRxuTiB9rMVPJqB3HNicrIXZ+Kw/1kPnej8q4+JI2QMBy+U
zDX/rBzDgtiE1ars4R+fxsUq8f/dzzQta2uD/DqFWYQx/hThEjZm4E5WmEQr5atC
sWgzyqmIkqgQL0Eh3iDrKy4pry+HFdLEBSiTdBT+uvb2CgWOR4PL/z3yHbnloKr6
oqQfvqvUOoc8hyJ03IZ29cKnVf1Zw14gYcRLiV97zIokZM753Vh3Ofh9ea0VkyzQ
sIlmX/P9T1WZzb8VGXLJPS2MFUxxkhP1gPrP7KPIVGdyTLhpqhxzpJ1waNVXHZq8
gPktAQBKc4eJ6RYmu1RQZoAVtq4Wk9fvwjfHu3B4sVw73P2vyhLDaTD3VyYQs+Vy
UR3zAdJgopHnpkUOCeRbkgsTCjLR/IwIQa8JFpJGOrAOdmRUwkFTO1tFawusjWWl
k6p1FWirhdvw22ylzcW4R1QLSj4B/FnWQB3RlLF0HzHSxYKOYQKeE64qj6pafzs0
rrOGoujm6pEGfO5Bu2O9IAF04lVBGjDIgA9aOaWMOMudjRb0U54Dsh8E/LbVeD8E
qMLbjWOoujW4vyQTxMG59cOnOPMfHdn2Et45bG9Ufbe+T/6IrSRtn7sDVZMFZqze
+OKcg+GCReInyLe8yXkxh7REuw8dHW4UFB0MPpbwuFj1AxEJsL+XbBW7OBMAVc1t
fRdsHDlUqZoGCaFr1TIjnf2oLKUF0ivBr194Cr9rTcmGAsALABbn7/hKh/JL+01h
lYpapiz9F9PiOwf2j+bq+r9u7G6DTizBGOWGRHEcxzsNPL9v424sDXjKa8RLHhaf
3o1HK0b3V9r5QW1pa9M0Lh9yAf9g/CPuS2L9wItc76ug4xZhVZI2rWkF3K4HPuCW
Sr6u9gO43bIGbvAE7LJ0Qaf167vfs4+cGSZZafqJe+28UbVBuSueuKttO5EhnM5b
BuDzvCpUf0NsrgoaubYE25KksCU/72Uj8xfZllAin6cZFUuqnF+D44jCtMg4joka
KoRRfnoe0RNjACiKT8HNQCjvKGq7XS0oUUQUfISgmE1ofVQ37NMMoMPNfaqX+2bd
pOquRVOgSyZFwA8qASnVPdLmTPWYN8G0K0kDmCQ0rrhLR7oyB7Fp9VZ/Vy5f2h8N
cKxtWHuFt4Kuf54PQODnz6BN3UwhzFtPjKZJK8W1rldDqVdXcVsXp9wAg3TyE2mX
Aewmt2yHlqWcqKN/IgHc9fvDIa8ZtfvkUyZHzhisYrdSgUaa0umgFnByx2V6o8vi
4CjbhsK/AWzNZGcRpx6W3HeweIuIQDK29iRk2fnrnvL7oBHNcOcU/wtxTWrsD7ZO
E+dd9h5/qohC//nupFyDaV6faZaaG1OUpQxvixGYPmqPBYYOJrS4IwSDbTpOmO+w
xRooQbgjbrzcrnKF7kTCbGgAMCJaB9dHOQOFzWCDD5I/FycHtbgNaiSYCbjcNvJT
KpXGgYzi5YipV/3RxfBAEIJQJYrulyWBshNReKIJ89q99sO3bm7TriiPO5sm/ycs
ogg0WG/rUvJfg+KgHKxfffRev0W8JUttt+CZAeX2MFfCK1UqFzdicPWd7y1adBGO
39HJV6Adwz1MAVnOgZUWw4RiHnbI1GPpaTXYsfALVamu0V85BK/IKNfU6n8YwJ4L
jd6q9R5mp8g6WCHlV9Cj4Dw1VGxUpBJ7wQ1pz6Rg/zmaxnkrqfueJXzrgaT2Kzrg
VX5bhoNgoqOL1S8Nh9bGRnleh7SiuvIj/lY+pDzw54ggm84GPqTIAfUhG0Al+G4Y
4i48OwWn0w0edlqw8md2RRvBe5zPXGTmsG3ARbL4lpd8Xbacmg2nw48iHKMejvzP
8BDSp2dcLemWw8qL0U4Y8EspLJ5M3QSKcKvJfT/Y+SrMgL9pRDJ8JA4vbGSW0avM
UWjVg5aqJDzkNnJCIK9++zZc2gVJh1APbMmFIXJNM/mccKkQdLp71mltCluq6Rj7
S+5938iV/oq1zUAUHzldp9feQGZPirVM4n8KhSGMc1+MnZm7CAel78zCa2kEkJc/
pk+iNQH/O/0erjLFIJotMeTIYzKe302+QbDGukfyC24Hd3H+kUXKGsSCnIptKT7I
0F/KJBgzeBykFqV6a7T5h0HalotjsnHSQ+Gp1SqV+iVmHYCaz4wcS/QVV+/lEsp9
oR3uiWJb3VlbrMkUHx8Fekud8ondEDpZI5sPfof1QvAbrM62r7HafGFxCMFS3qjD
ObZGAtUFlucIaIOYSmhtDsUr5KlR5LyWOy8i/bi3qj6RoinEHmy6AzZvWxwqmmbS
SzkmYOJPRQAWTP7Nlxzmg6nz+3IuGPwo3tCQF+nu+C6uSRuqb+qmX+roUMy8Dnx5
pHmEA2mbPnL5gWtpPhh+bfFwD1R7mdYKeNcLLcEn6ezLcLvHTPy632cOvOabxDHJ
9e6J8J1mg5qFP7xhCjdym4V3oHaPufzb4B8V5lvNMmIGuWpS8q2iTxBcUpUAhzLT
SCHOQPzudlqgo8Q2+EtXq0vkPDIHpqja442CgRATcJfo7s9rgAEfXVCQ5J+gBYsz
arELGmRytqOcayxT1fKOI9ubUwP9DFzvaeFcxJbNMIPx1x2hHsQ6U7mE2pgqNF+x
JzwvXLd65fQLkyblbWNjDc8wqAZHoNXe4vNT2MOYh2noVMatHmeZPPUTC1KeGpsL
LrEdBa8N4UOqORXdt7zHGm6iiswAp3YnRkgbeUwoRy7/Taaxtkfhtfdvhgz1QZEa
vskEYqOMT8k4WMsPm7C6IXnLg6XEY0gX/4egS0G63tpMX2z0PcjsTUXYM4qfrNEJ
t83VLjRcSNDD2TqFvb1vAN1Eta4APTHPmmBEI+k3M5msb2s05pccS66RnasuA9Yy
ngIZ8udO6g87ixzIrBAB7GZCwkforyPlNZOwhwjO67lFg4xUaiD47/v+bjNOHiOj
sbKR7PcBogjC+zQ6dNiE2zu7GGlLQQkXmWqpqcN7XNPE/zpLMOpxQCwEfzPSFTxE
pQBG6QCg4KaLmGLnd2dCsseAM+O45cG46GxglmVNX1ekhKl/uhf2a0tH/tasgA9t
G2QM5AHjfeorROPM5KSaAoyTWu7lA4Oe+Z9hBJEA1NGtuI55iP/3yT9nDM215pvM
oGwak8doYw4Ia8oXjb/J51BH5+uFgUKZ/VeFvN5W/EBr7gLIfAFUj/0aKZiQJe/V
eIaPbNzDs1Srz/HtNZ3YraB+ApTG7yBaLVkU/rocwUjfTGDHipzVlB97n8iVo07D
RnDLefs1e7qAY+CPRz4zFgoAilqlOp46RJJZzJSDxEaRyEHGWxoF7EAdR41X/9Pj
UXUA4YrCuUTLFbPj0Bg7xzVIef4FlgFEu6+3dfKCaaAthagYyf2NKXYn4vtgVUZl
NeKeowvMM2GdXdU//a1YtuxRrwXUBW0FawK0IgdWDK+cXnh2aQ5DY0WcWCZxQ63b
cRScave19/Qah4e3aM1HmQz1zp2+hDJkQlrb0OOAN4wYPJUxrIXRepfRftUkQ7xb
w2QCJmywKfzwOIjEmRGtJsrN+yGzhDd39o6RWC0JX+K38Xs1lFTuvvv6B19dZ5PO
xw9RkozzvPBhaPgb01YYvz6+9NttKf9zmWSXjPV3i/0KLmDNDxeFncIsKoj3PdG4
gj/fC0qMr0Obx8+NEnU8/v48cF8tYMjPNAq8ZhaFqsGVnt52Dcn3ssxaLF0AeDSQ
JwV6CeiqVdqmfZJ4fKac3YVbA9TRJ/LMre4FiE2LCXfYEz+k/SFWm3Uo1yr5Q7W5
5CeTrusPpd4oXzgxyvRI2/BvUQGXprRcFo+n9T1ij+QbbX7DqFiuoxuwRswLrqa3
UvhLdcZuXlHpdNIIT/EX+fea8aUt6h560xZrQscVFI3/a5ss/l9PtqBQXiIM0zOI
C1MqWjR8VRWDrNj3CpR01uaM4AB7D9jHUKVue/lfXC1nPihT5M4owL4H8GMAmPVc
oLh6BCM9wdEpjHYW7G+0JL7DuZW7Ldckf8ifi2e+mCpGmEo2CU65dBd/H5/nAvo0
B3zHerJY/2Bh1rdZjiGEIAOD35Qm4AdCE4XxqUgYWvdjxx8g3sg7MBjwuoc9x8gE
BNwitznfm4dM3cCoUvrPUjVWpOcwQD2UjK5e0xDQcVSfKr8TTviZNYanxm+jU4i+
KK1iIfZ64ZS2qGymP76mA4O1Juj3fHFp3br8PeU4Mzff9lT5eNZJZPA4/IQUWX2U
wZNjXdS8T8yjP33K5dIIEFuRW+GyJUEs3RPaLwwpMp2e/4CJ6/Owq3+U3yo2OwBR
lOo+xUtMhRtbQCke5X52zgjCa0JQiFT8SZC8GziWA/anpqn40Ze+O1BEGRludYuw
dfVZqfa+1HnE6n9KTK0qFVqxM925GGzVV/eWTCVjKIIfxhBuhAImcgYKG8LL5WHa
G5wDJR6NLQTV9mrz50okO8vlaL24IF2muUNzUAC+TMvVucajOVp8Ol3etC3VgnNx
pKRLF2hyW/sr7zm1RNqRB2GEQ/1b9hT+gGfsBcxsS6vpPmrx7/4iB7CT9apVcIYK
iYnTEXridnaaHevYd5uRFSv2NiCjOmcoWUBac5idb7gZOZzB7auxn+C9Lrn2NqIA
z3+OnLSW3PiU2EQD+2B1DTwyY3vM8zalLcJ9uJiEJnEmAWBLsUEESkwVS2TGAtnb
/vH4QfY7DYN5uN618gSFftTrZG04x2LCX/b0WRfe8QZZLywao+5N6EZfFHkKF90Q
XwlS+hGEirKMoOg231SUoHNwf+x3Z/oeWhz1j+WlStX3q5O8kv9XQhf07h2U5YuL
mqjj0MJW6fvKzZaFwGEU8cPEP/7SAHvteUti8xYVEuVHkY+ubm1ar5joy/9nYMph
qyTdzO95ojMd9KL12u6YMk9bO/ny2mrUmzJYPy9BR/obRepjiuwG8CU5Ca8x1HQU
csQRC5jZOKJDWmvDHFVC/hyf81ESKMYidx1bo22l21mbw6QAj4qK0JITPOzjwI+m
fojr+A8451cvMUkcjofz40QxG6uZ2qJjS5HnYQRpElJZLpL+ZX49VNyh5DyKGACf
zlcGZz+Nj85dMpvjVjuFtsKvIHfKo/zV6uo1UzRkORT+9WeM0fHzupDmqPme16Jb
i16/aTnCCnOJnMadIuj7wl7ZOB8N+IeLpqSmHQC/3eBDTg5ihCWUl2J3K2YhgMm7
UDh2vp8oymRF0un1aWamBXO7kekHr4E8/gz60VFnLfbQEzoA3OS2Upkyg1HK1t+w
MWLY/ibKC+nqoDUuzV29mspculQb46DbSVc0UMf35SuC/ITLLdfsmDXyqc31IViC
ihaCez/DLZ4aDOg11bcyppyKJdT5ZJZOVL8VzIQ1g6ZjOlyM97Y4MdFEoFdfH6E3
oikClIMUTedHtK19wdq6svwxiwgqTRD0CQBtF8Glqoppqyy7/LhT/5x2Cmq08vh3
bPrCue6OeSBmWBHeUJM/GJaYxFEqzdm2Rq5Lgn/irbWIY6qBRsDLL6MsxLJLoKoQ
t4kMUL50PtTYvg48LxVy6T83N5ywy1daVaz9HTW6U3uKw4UigR7GD7VGUhbA7wta
X/jMY7enUKui4fo/fth+5JPJHgh9O1ZUebR6SPsxNIgKiwYCu3ShEEBFTnzKT95+
gtf/FpngvXs12n20VtQX8+sabUtKuzD+MdkawKJEAT1d8zfk35LFKu9Fw1nsT0+w
zyHpWt7BQ8ALG56q7sW/MVm7sdpwnv5xrVQblazTcAGtn5sukmqot+kr8k1NBdj/
rzxborJEYePdyoWLVawy+cAvZnBXdioFxlVLGzXkEhk07LG3nLu9m+ZY8Li5StH+
ztoMdNO7ODgAacBORi7j3GeuOquEKaNdMmEJ4CdAUJvoMaDWW55Uqpy44rE4Snun
7IC3hw/HvUCs4e9d4QAMLq+ee0nNDlZtha1swxgUiFfStzD++GuErZnhdUhkz/f8
f0sAkVxqnmmzircdbuxXq+DdXe2g0/hV9xglAaCmF2N01XPx0Yyo4WQzA4HzZXz3
Up9COPeO4cJMLur0NYyLp7hmuajLSSC55r3DLCznPzI/bz1jpuTSg/WE+mZxM+oh
WlmrdfrLej1CrhjygaFlUsSNaDR1D4hYgtKxO0vDlezo2+1ZB8MVjWDS9pBN3/0T
DCvSKeXzJI9UGEMq2Hl4W8a/PCDutWgs2ZNub6f/QjLrWBwPGdiBTQ9D+lc9JcbA
6RTX3Czeg9tNp9jCJy9xiEOix8b4Vv8tYYsbNxI+HaScg1Lyx+a3DzRU94aJSt+m
FrZEPV4/EM+qi8SCv5yiulBhlfQPl7m3YOWtuYz6AzYR/xqTQucMI552m8COTiYL
Ok8aQXFztrGXxYPON8yQpzuB0Ry1gJDP66E6OviYqWLUuAfj5aF24jqe4XgIE9n4
Qd7u5aJa012YC+3b3oHV2yJJaO0yth6vD+riSTPT16GF9brRrPShSph1UlUTKOnq
L4fl4rvqQJYlmI19zUl+GrhQKVohDt5/4A1vJCDbgmp0XnfZdNOWHErjUBfWEavU
BBam1KTwAsiknJSQK7Y/IpogHal9/SmaurBaFzHZBBGyAHIi1+/+anjieN/0zoaG
Cgg2tCf9yuIgq0U7/N+4AERttWB1j1EIeSjNzPcaCVOSHLVLsm3ax8uRkl+urc2f
m23hdBHGgPwhziSGpkI0WJ0Y0oeI5a9pBQT3B95k+uHEQ9o7KThLPFCS8sfwnwPk
o7FjozQJfhIP3YMO9WZYvxA7Avqew6F2iYaOKxlcldMKVMXCO//NQKuy4N+Ymzde
r7LyA5x5mUvKhDR+vnBoJvO0Urrx+JSlQfk1Fns6fC0ODmj8B5MbBD0mDZDQqxFf
t/eI6KbL6XWawFTt/5TuJBkk/su0Q1PuM19gLNT81VUl0jlu7CFqLbsaI/BLzgpw
iDNDIEPUkiNdzANEkfuhaNOok3bdmarRPEdvV+YyqhZcne6HxE5jN5dVNQihL/0D
+VyIUdXTLo1A7TrHruznV2SCEOJYe/yv0rPG8at7uv8Sa6W0fTQ4jG+f5vMT0OgZ
84wEQc1y0v3E80pDtBBNfYn3oceDm1hcbINM4lcjkFErfHyRwok523f2Mr1aMjLb
WCFeWZBlS+HpfNL/aIvVZJPVJWLfce1zkkoJRABenfdForbStjm9RDfZ0Tn/pUmx
Npwy2BJt5BW0cS3oQF6yURHTBsIkDXmMQY1OjJVZYpzPdB5CZelYDkmmMp4h7Z9D
Rp0t8Azn1j9mKLXV0Em/vV2FN1uE/EEV0lECjkxqs/yxFkjLd2D4+7ewHFeqWoRy
RErUjNBv5Vj2rHqBNdRFXAyafCbv5u4GTilELm1v9pEEW/kRvSCNEU1hZ63Ajo1P
4mQ61tbZA2RewIQ9LlPMqAGvCg7VrN/u3fTHG5P4kt1spOaFSbXQVHasHXqurFNZ
Jua+ugyQwxBFjn8yEJGeIt4qTdG36FrHf+dlLO8M3gD/prxVQ2CwsDfWWe0hCiVy
s8fBMP5z9UkF0zBKyHP6bmErIRFkLYukdaoSdWcpdsrzw4f3ZbSFTE0wW/3tyRl9
JWKlEobG0BlCKdLeT5QQ/D9yQrqgPxAPhYVHY6EoFEYQN8SRsHkH818EWwpRt3c4
naLAwTOs8925Rl2vGHsW87qaSGCod8PmCHe0bwOgzexJZqq4Z7q4FPoXVekSBDkf
rfs4C/TvGBb5sMo8ZLRzVfvzrGo0LvbOEAoOrWCMWFxnqYVSlCTd3s6J6v/fb27I
omeyNpAFMpZa1RLizBD9sZAqDDae7WHtxGshHmdFT2JHSFkIOrV+XVdubrfV6m4B
ngt/rM4y3LGFORhA7ZQNxAwNRY+40kZWSQdW8xjh+N+zyYKoYYcqml3S7Wtmz6US
xmmCEav7+ExGJSiWKaC9fnT1lrIib2CyBTlYrkRN7nPoU+7/5qHUIQizueFZzRLF
l0w8mNH/HARNY98SEY9Q3+ZeumEqAcBevo0s/ohtz33XE9YMp2PdH1ih96/1xwwd
GoYRXeWVTKpi7Imrj00CZLpsOvZjr0roC3MZU6dhSq9J9AOc1AB6zdJY1QEm71FP
u3yp1csZlIO6L1miFkZjmmoUsRyC62bz7IPNIZDJam2npwf24YHp0x2rvpJ6yN8n
BcgQUtUfxGjkcgOO3MnZQVgC3MmDJdIMaVjE1bFqwF+sbuGJUHNveNyYtXJ/AFQ4
WwYlqOoy5CpD7ILv24pjKVTIa2/gtNjlBBy3hNGTop56zM3Fj4Mj9ByVk0GqQzRS
YKmGL52/ZHoRqZwM0lXTLmrgL4axiaYtRhv++WBOk3EA7g2oj792V2NvVQJ/YUgH
vX0Sg7jUnr5HYLq5FVTj4MYo9GxEKDxGXSAAmJlvKQvvPQyB6OrLJbYu/PS+S7DQ
NofZJ8+KwVgr0drLOPofbuar0DVMLCFVwVEWpTEIoJmxuCDtB8jgnCLatYYQ+Y3L
H0ikrDtt/NYx6g2E5JYlxnYjbX1aqa3LzpEA97LUdaYOZ30AksbMfAbqbBd5peaI
DLJgtoglThJMKwu6lzOUW3RmyY6uJ/uSQWNSPzT9jSTIN4s8w+onsXZ0o47xEkxA
l/LYOQM4ICVRpYv+XEAITnG939pun0JwpgdQ+fEHyR4dORui1HXPL0cmxjgGqmyB
W6jckQZ+J4yzGrvHOExleMD2SRyqajxNpP8+GZuma5gIRyuxazCioWzJ6QiewVOg
DzP5N3r2frXMfn7DfuD6TyTcAZron854sQ1Ncs4HYtMSZ/8qtVb1x2XhCjWm4Kmw
iCc9kdAzR2E1Gg7wcoJdG3EBJxxaUAepP7cFSywMAkWcTUssGyF/4tqgloR5jwsO
/ZnPucwZiWJSOAgjY6Mni01iVGJ0hFhLILJqeltKzZzPqeyWO+yRPgPdTD2D65n3
03TtBequ4usZhcNUfnDLeHZbqOq6WHhip3p/azrCo0MrLQjjVx/NzlWhjw/Ho6/D
Mzspn2bjVXl5OYkZ8c7BrRUWA06VCQQ2xkIjzKv0PlVeRZCvtLt2NeEtMvqrXRiS
GQJsambvjMPoEH9PgRQ7yn33AKqqqcS3CpLCEN3T1dZx6bBO1xStnYLkO77thGZW
kZ8NelLcK+4RH98MjZdNagGAaWs8K5pO2eUpF5WVJnLAm2TxTIcvq6c4XdT8CvlZ
Dujk0bDgny1ELpyWeXUDtoJ6JbCcYUyfgnqTB5aVJrTDyuHImOLCN4zfg+Nr1TXE
VBl1k5x1JD5QNvs6n3m8hyz2iOyN1QtxBUayNLc+D5yK8aplkTOhr7Cp7TdJkfqL
eazUp3wk2oOAfQydjRX6dzvmxxfaj8Jd9GJi/0N0fon9W5gkj/n2qb+Om78ye9OF
aDrglsuUoL0HVXrH8l9I3H7yztrSM/xLVihy7Wpa1+VHl5v0hx9BGrzu+i+Amiao
D1cFs+i1HAVv4kBpJ3cRWGtbapAWwrTKFg36lJ5gM4qlOynHOJ2FM9e0WrMVl8bi
gRZ8TJcrMefx4U6XZ7ZUWY95Ygxre+nR7KZUfhNMcdsQrkB6JkbXZslfcpzJuP8f
9M+818AnRjiQYtR4KFZOETW1a5RsWFyVq4vBXTYpkNb+1yjFj/DucHRwZWubBnuc
lv4cdTBqXT1PxVV4gbQE/LyxcR14ScXmDGiFhdUK6zPD7rk7QZsBK9jzZ7+DGY+n
SvVjs43U9eBBZF7HVivKqZjnIAtFmecn9+YgR6AOE+FOg4cWr1AXYATePIdmlUVj
dk7C0BbwArHmW8Ffw152QdD4SolaGEAjvkZbq+KTjV6MeqyS572ppraDDtGulvoj
CmMbjTA/dwasZVS9APTCdqGzduNCa9kWtydNBiEs42qjGM294ttLagzzispDep5Y
jzOpBQ9UUqAyBckyd1OUCwwciteMAvFRRx2WbSXrzL5fzznPqTv0A505ruIMKyf4
S1kK0rBlPG+bpvNkPsJ1Pm2mOSVaDxxqI89URi8PjuvSZzGn3z7cGgYusvybJStZ
CKDfv8C4vPAOpsfKytmDdATprFY7CJh4zw0VlWBiL43HOM6BA/HjtN2cvDM0ZOoH
5HBSNoHwXs4ftiYbBtfLIt2kRVq/wvBrZrfO6YdlJqlBEVSgkHvxZiBh9sVtqB1+
Q87ybU6biXrMj8H67JTPl27J5So/OKnDGyaFFMfN9Nb8g1jExSxnVQ4lH+0WcKbS
/kfZqvG2xyOyo1OFANUmc1IUczH+HBRNVOJwsGk/mv/aJVnyYj8aLozGL7xR+Hg6
LSV41uwFpmHEhxlbeBO3EXWWl6zin4fnsGlP/pNgVV7CGeNfuFqMUGjyIAJS7sMR
Duaq59PCU9xdjomias0OfyC5QN37J5SJ1SApxfpq0lRmY8+yXzrk52oj/3PQBbMs
/9UkDwzcCSM6miBOJojUhACZCDBc3B/AH5J+uxejIE6JxtjGZ2wzMT8tXK0zIea9
pvxzVIW4yWLlht/LIOk91/3rEQtVgGJEISEXDFQS/ykkfIYvAyvGmwO8tQJbgBdw
kXMpE3DQIjtop+8NajgR+rGFXR5HTDqapBtuKAf6DdodrYDMGEaZXm+u0q1Xbjhp
QrMPJCuSXxicwomWX+9KwQ/6KbtUf85I7/7BfvpGEZiozIYykCvh/2oIJI7TF1pf
44NdFZOJT0VxNkrtZbDDsNOz3KMb5J50JZ3JfRTp+o4Vc1mxEe/ePY07sI7ItN+S
xFllHaF4A6Rjp73RsbKWy6CZ56oDHQrLGsUqSjr4ismqM0YlONqS3fCIcOv2HkKL
4W7QReaneflh2drqnjaB8wnIiig/0SPwPPkf4IQo0SRVOup1Pz8t6gMoRTtcfAJP
XBGpcyhZ7Lz8ipWPBgOowItnDg612u9dVDqDQUIjUx6UG78rai3Y5YPoyAh2OTa7
BDiYOzJA77KUSijdRvt90XrfxN6Fx4tWcmmwuN1miN2lyz5KQxNTDbNbfsxrKFjj
rAjxKPwpXjrpFAtAmfS1lSOjxfsmzPdSfQmm4M/qhsPHfHxpm2ZHHpdmlXs3MGs4
Ki3hEdTT3xTBNE/e5j7ykQL9lizN8NmeqGZy7rl5ft600NG+9HaCH7wzJSCGTIAE
zzkEXuuTnxfG6Rfalk0jgDuASsSSazvu2FGAkmvvhunt2meApRH1AG52SWTEZPwE
hQxcERvVxzJjfayZm9yT/cNwnAtcHC5EiVBgLjz5upipNEezvsAzjTDJmZbfyIYK
qFflP6BWxPt4pIMNdrwb+Jk3jcTURGAbsSsNyvqAiob2Hs5ulGENg/syXN8x3XWJ
zdrjfgGPn6KZtHU5S6CL0NKkgH1zXHheD7AA2Uic8+OZf75VbHpMb3uwV6fQMQQR
0KC3kn+sjoyHeYyIKl636wdUsNMF+4Gr6Zc5Q/fhhK7VtT7s8GK98E+yTY68+RV9
m83HgM5iRNP7jAwUQTojKXCMJjJIhaQCZz4+7ObJAcahJCULp+9whqGJ3DANa9iE
OO+b2rLL/uZ1Xaek9WqmMzxj+MDxax/8qyyJTx61Y23ErQqhyjFnzwm/jOrigxmt
29VMYFlrQcQRxxp+Wl2iMFJvRpmIOK8D4xCeD0Mh+PRZaMLq7fFl6703Gse6nxsK
03Mt+qatqUd+7DKR/vM+gLSuS9dIIoquKnGjxHtXU7umheXFBxot4AhKRyCFsaU/
PNfNiC/HQQuCuODWLJtjaVSCVWbfW6W4inD4wvacb4wIj61VL/uwVmxMelNxmmYt
BXa1KlPo7kwHLbY9H6s1l5nfyjE8/RNi2//+yy2bW2GQMIKUq68GR6YyEthgiefb
e5S9ehjoKad9ShGZCiuvZVQ02xteazLEpaKsc36kAC6tTc5z6y12uyGP3sqY3LG1
6/NbOtBMpTLUogjHGm0/KWt+RYlLV+ViLt2YLXkE6F3Vx7rn1nQvvGM89o293bzx
yswYcbexfmHVWa/ngcJlZBAW+uUECeF+idjwCh60xgLk37gZU624fWNXuC7AG4lB
aG2jgohr6ryWNzfHi9K4Mu851+FXkTqidU6ZtiXuzgIkcNYZKa7FVb+Fb91uDh8h
KxV055mFAr4O4TdV1C60EXTdfPaclyrm93QqtRlN1hN8qXPKrHH2Bo9yKOVBvWXU
jHZO/6sGx2tlJuwk9XOHPo/JyN2Wtb01+Ks+6Jle9itYkB5/xCSuA+XAT7ogMnhJ
xnjMJMEFeZBjMnzbpYO8zBoaiOKsP64oGTOnsdsQNLBTlhsx3ecyozdf9sQgHqsF
jUStzfgy013VDwHrZhx5wXPDlr7hkxUxnfSpcB6FaSeVlAW0DVj/BXM+P+neAUDw
HubgR282kN+aeSBlFEfutD6h+rrA8pE3V6rp7ymF0LjVEE5PjIKwZYW2QO5a1tD/
1c1Fe2+JPKjPx5Rm1mc+3Mvp/Fj6IyCkba/6jgtE5n2BMDK8GYoRE7GJjQxM3lLY
IsJlLjEcqfHLYHJEG1Xb4glx8p96bfIFYGFgpoeObq/xBCesJkpuhbFdQB14KVGw
tPsJU313oG5pZvPWiU0pva4qwUTUiP0+SjMXOjGPHPD7rkm2/XzjHs48YqI9Tvr8
Bi0e0Ubtsu1IuFrETddySwwthvDEZ9l2DjhKSbJ/RYUMtgyU9X3qS3Lky9NvTfee
CAKGw53IHvrI6OztFgvIDUFvxfe6h+E+UoKHhEQDGSuA/pyd84G84gBQC5a7/0Fm
LKW8VU7HdsjvFRxCKWRbW8o2WsGqET7VyJfhCvg1zFAKKvZzvR4GLyVxxKNCzWds
FM3byPFaQasQJg7HvaQ13RXYVbcvK+Z35golPKBhBDOqL1fUN5NT3sVyANZT1osi
l9svbPM9Koj0IWi8eJ9uhEL7ZHSp/dy+OEgrCnCDnTwyx6qH7MLRvbNNbBAQze7J
dWW1Vp2M2A5VUs1IQrjtMc30oJcdS74Z50JCYxRnCBSt73pJCM1Ttebi5tvV657j
4WWQZbVCu2ynDcReLQq3TJ1fS6YKJORfPNpyM0N57HyG4Ztxd2uJQjVuqDibUTlc
mU/r8j2tnbPatYWRUaBU5bVMcR+LlnFY3GXv8A3eKJcFuxMu8t47C57c750srU8i
QwPGHvQVigtpc8DCyDGk4oko/AhZk8jFTtRbgkD/uFXhyVG6PNcomnYSkcdN7t1y
QMb4fe1EGOC1krQlxROFiPuTe/0NQVQ1z7GFxFeWhwOHIPkA2Rdd0wXt0vCm0iPp
z/3xgD3d+k57A/wgCkaX/EWKO3+SUL0Q2it6N5NGlE2MseLTF2cuiK2FflghqyX/
TDG6GMWjnWxk2RM2p1IWMUubiF3ThdiLj0Mt0nb4qPCBxXcKAPps4gJ/OMVR4z1C
PsXYbWsH0hdQqWiNmbR2FF8AnADiJxCYDbWVir+CGudrry+G2u7etRuGsibwUmbQ
1QS1JrE1yvQjHBJlGwz7pBEzFHvwjQ5Vomd+Iji1+dpb61gaDtj2vwTQkHpImJn+
pLiNjIYM4BoD3yICh6hEIQkqzWCMqPs+Cy3hKWk9xMIvd73A3YmVKnztHF2AvVvR
GZiPIJ36NZ/9mO5g/FwwSaSNfFTXvAL18MUMnei5rF2oPAgL1GPUXP+gqURB3DKW
Yq3ElVDmUs8Ce47t5lXlA811EwZnBQEk6Tt59/5TJa67r842GsQfjdNZaltQHZll
Ga6wOcvBHlNUsylTTiLT+iKDZ06v+eI7VLda4JrHEJiUEcnjeQovTXg/4X3EM2ld
eqn44324xMjoHpQlT9sa6D7PXIC2FMilH9PEULmigvVMBepy/NCipgbo/f3ny0lD
ohgHy3WVHsurC+SX2Lsdg+9w4HOTUP5PBMA6PC0UsBWaBsPpWF+b2aQkm0McCwi5
hdObgQ1UeoydptVXimqJteqYBnEQRjQuSrIwkGsCp60kwhA7CYV58kyYnY14443m
/5lPjmlSWVk/MPFI4NQ+FQWXGm3NGHXUGPbvUtoyxDjmKZkA44bb9qcDTxHVqKA6
4mlL/Yp0G6RQV0/DRAW4Wq6PjcySlIGDIN2Kbjr0AFtjLXiKu+Aa5uy1fUM8SKUE
eNx7sUoIosVC5LlkSzBc1nxcIhotakRNg45Mv9jGBqXgjnEcIyzwP3JuGdju5k88
WVyctKfdJ13RoS5nHsp/hPQl3F/vudBBB0PePQbesNtky9CIeju2FMMAiqQsaUoz
06GFeXozsiGZBdmP1b0cZGnL478Q5eJfgxZJ0NKV/1nyudlDSy9ymN94mudj1PNX
OYjDCVaOgBMZIEVxjblQJkMltadPfPA8Hf4V+poe1eB9mDb39bafbVTxEHCgBG8s
BwBEz1ApxT0j2FzrPAU3rw9dAo/ZHIVIY+nLC+rdkCXL5Enje5VpqdHraoa06Cxi
v4u8rRTfTCPz/cx9gb1H67FV4WnsEedjOufaojJCtdJEPn7S3T7yaNJ7Q8sPhcjP
tS+1/rTCWDHAjMjH/ydWWvCuhf+3//kcqAxA8NyjmVTv9exQIz3ppG1WsfL2q6ig
7mlTooPGyAYLGG9eVcIN0V8YIp8++W8svtf+qq9I8GmOg+ii7SRztABO3JDw/L6f
RudLvLHBNCwf+cfyfmx2xqXcVwa6IK40Js3/YbGO+E32MYW2zNDNbCqJ10Oott+a
mREelTTYlnaK7LDBjKvs98ImPJlDC4662NnlehnWxcY7XTZm5VlndorFkvoLFFWE
BOUpPFZkss2lKM4eJGJWZitVIe1ni2MujgaBgN3Eg3JGY87cfLIdyQalh90DcrLb
rzbXt6wW1isR7/7YqmHkwUsVJuZto6Iy0fidoGQXgZIb8kll0Z2HGRNfpkCifcg/
a3UrKS+TZxuVlCOmMsNcrXeiziQmfqhyi/u65l+05YGIUXKxk6B9RxfDBkFlbn63
FaD5izAiWa3bxGkKycOpoi/H3GFYTPbBDi8NQfhKrYzYHdSpSRjm+imQIRfDHD98
MU7cnsa9Ol5xwcWs01ISrFdEQW0OwwgOnjmd6a4ZbpcAh6iOCwuKX1nKiL3WrEIS
oD3H0oPWnuO8EhX7XWyxDgpTWRyJhDhvSBVdrduHy1gP2tPH7yqMxHYxkmpvffaV
/fTaYA51DYxYelWVVGzX71euLzoPgDaHp0wvAiyKttUU6cwQFBuRGOhHGYofPm7T
Zxux23CnhAsmyooTpGe0MVA4FxA6QrGZ4CAzbnUCibG7c+5O1CpAeKWc19o7kQnc
8MmDm8+CIk6TwY8F/iBYm+QnR1VT5uQV1Sh86OiWorGOxmyGu5gDDgwC77QfeZGg
m2LxoX88WKP3qBLZ2hpQHQZWDsBYLNWReVQkvzCS46MIeSNKOTD8tTIXRTQH2bj/
GXKvhqe39gx5iErkfP8iMqUaOWkTBuUXzOCFkfXWjdfclu/Mo9MoWanapZsZE8jH
ywXLIiUV0fj3Hjs+awlENQXMyQ6I9tYI2Gw+5n1ZaV0CjnFCkXA+hm+CVH2wTZBJ
eEwMy2J/evaVemO2J5aVpPrZ28gUqBvgUP73Wh/nO/jF4tdbQlN322t2qZo3fFnm
1+jDAW+4tKc+mZRrPYFWbVvawcu9x8qYYk4ZSlGyIg386yd9Agtm/9Vk18lK9nmw
SQLTaSLPMailkkcmekwfbLnt7qY1NrTTLpl7QlPDPB3WrpqgtRf3vMi181CHN0+R
f+k05PnwYol9i8XYzk8juBJ3ts8uGeC5kr06mxFtm2+L79nwRYQIw/I2Aa8qJV84
kwRQp20kO9LE5zqZTSA3Vq013IH7vqTTJqXXiE8orzY5So8923l10uKH5EsTuHm2
tx6qeW2WfV51zAjItb4zym93MiKFjk6mdNFCYwPka8hs+0Y0QzBOBYEpcGDsIDaB
WJnmUKN4Ry9mFuMqQr8L0qJQBapLewus+qW0tMfb/N1XINABijPDrzKfdTQqerN4
qo2jTjMCAwu4v1QfHTa0VbRxQE+xJx3D9y9JPVZhAfwyuMRJqHzKjgh08/iX3Klj
Ltno1kIpaMIy7UKYjgmrKzM7f8NfNRKDSBdJ87I7vSs=
`pragma protect end_protected
