// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:38 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EbngFsVekMv5SUaKgaM0HeG3qMLE3L4Srx0dHgMFvi7qFsszDeFzX0LeH0duoezn
ScTOcWokO1Per+gYqApxUWEKa8UiDgD4PuhrMpzyegS9boTF62S+UrE9wKymfkVi
a5uUnD3DcFHX+8vWSezqR2mzPlQGRJhidzJ4orsxm/U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7712)
rFf7d2mGKzU0TNvIIMApiBaujs7TamRKqH9ye6pR+bVIp1HA1lijvOuTENUB5qz6
fJ3k9MAtJ3b5fV1p/Q1Obg4SRmFvlDD/zgx3lnozblWapZySFRYS/OLN/4h8loL+
Hct87fywUfkoyK6cR3HrhflMVZIsfq4hjopwKNBa/7ky1yLzAF1QjNdQjwjKeF9X
ejqiQabmHn6wdDAru1TacDjN3Ml69tGLpl29KCSE18vz5vgHJ4hPDkfEvG3jXWev
FkwgSqLkfGyaRTLnNofJe+09lofX2v/z/eTJ6FQk9tpUpaXEZ3/gNDGpkdZJTLkz
2E48h3JsVVksDMVjGb7+7E+65stEh7JW+iGNcaLS2wZCWothyNe4k0lBuAnEsaEp
uZttrjnspnud6/SFmmt2AwGXA/ucaRvPQ4zHfTLMhBQIPhzG9XWbawYQm6o47e6Z
pom5TlDqzLzfdR0RHTUoKum/nXc29HTgJuRdxH1hy5B8jikF/+4WVfPG8jaoXHNh
RXPR8VOTVUqHu/cWG5yKdeZ8V534dWrV2PcSJL01Y4iKBsdcjuylJKOL70XzHmu1
B7UOSUugmEP6eD3PIBi00a/RBZ9K4oD2pQNR5ibc3q1oRywHACBCS77ndYhlvwB/
8jHIGeUpeljIJVQLb+VS16mZyRqCvWUQRnnuCmjUch04zhdy3WvrnVwOgYEw7edh
zWxSAZgFvMun9CTGduQW+cZXGYnwo/e90DUcbNgH7bjHEnFv6F43OFzGBXU8wTzn
qi0uXqygOSthv113VzGBOAnymsJVhjj2lXjUiTD0js4B4a/m5KhoNsS1bMCiCi3+
uAxdfww3EBifngkysVen+U4TDeRb1MylY1gBz87PZ5M0csTHulOMew20W9z496+r
vX0jO9CSxTD9xlZYm/+Niuzizk2/f+9kaOENWAmxjjbMEUvd6TOVZdj0qaIZOK9f
Dj0rTre/3oS4IoE0MqEUCr6u7LA0UvnjM2uJfLc1LWv0Y2kG6dobqTcnXjftEH/5
y3vARlw2V/fdMtYnX7G5wgE7F2Q5DIcPW1tSrB+NOyZrkXsvNdzHUifC/p/+9wfP
85NFlc+fMIPwx4XeViCBW5TWNdgApyqvli9GpcAwSvIkpRglj6aWejh2U3N1DqzG
yHtqp8f05YQKyh+7M0asq9/Q2ORl03RIkAgyN7qAfdpOh+K++UAI+NGudBV98VeZ
uC7RodQjGN6Sduj7MXuMcfeqSfW1owErFm65VjzE5EXHGzO1FH0p4Mwho0Kc3vNw
YxQeyy6M6JMv374O8wIUKTMqC+k+FhG1RZXKlHuPheHRO25WGhfQKo0ORFsW/gFo
eANkPKyzpwZ+y0m+IDq/0cZccL8WOHsTaf5w1OOm+oO/O+shvsItqtjjPO83oIFE
JcadDVT+ZK5FGNYvxRGNeQIF525uHp77IFO7V+B/0/CoCf1S61jaxeW6WZjzrucy
qcjJ4nLke0cklXYuADBgWrUy9/a3xy+sfblmaVFsKrr+MyKgYtomUG5r+K9awB5Z
lKE5preXjgDD6+5I7QYsWmDyq3v6lAriD2GKhqi1au5MMkV55SemzrTJu3dCIPRN
yiMaBiZq+gxsKwIHyP5stOkKfS9DYWpuOvyekFbfYhv7ZxlAFFSkIxLxp6idmsNT
SujsWdSZVWaBlXQr7QANMy2stY9IEOT3KGjBQVki+PA0DEcQdp66XLtE/ur9io/f
vWN0MdwIbZT0Mzn99M/9rCJkjJzS6jAD2zfL8HwVuajx9OS39ZK+EJ+m3KTJuMl8
9IbhswmNaa0RyFNTaMcEHA1bxLl7lSMcG7XZpC9NJVQzOXaGmv78n7UO6yLWMUhh
wYZunZIStjmI7iY89XMI01o/vNTTMTvHrZL6BSj8Zl3MIyGxW0qgg3MMs9u2+gq+
qWkA5OngQjSMLP+B41LtwXpaCN5ySiaYpxRKU5VtQ9dfPscdkKbrHlGi72sUce+J
QZa3cNkOFYpL9TkTHpdRDsFqvtJ2TAEy1qFXoLwYfq8eXsqZQ4KHDvtL1dHb2qas
1H1nmltFwY3YqG1mZVmc4I9rLdBX23xLNBWgTIs/cEGokE1KlPNDasaGyvUdG4L7
nOH8rL7Tq5GGKNLQ3AQTi6VKY3yUQ8f3cwKdkya1d0+LdIaxnl9UixIfjwhsN2YE
ky2p0Zs1kl4991kgmx55MZyNzGLCwQiathdvoOwsyGkR436CWdVj93Lpgga679ax
HNJbl0vtIGoQaOailPVGqd2F6xKdPDuuhf++x/tsZbv3bGP5zEbSHxHxaK63YfgS
FxdHXj69XRw6hDGZdATNTU5S/nQ7mEp4rvosNldnmKvGJaf9OcQFtl2/rM02u3E/
poqmVxjkdwhYiMnUuvH5krT0OdG0X1BPUl8cXbMs8BU7YU3SkEy28MdYq1vKcNb7
SDyBb+tETqqb1u/NwaKd2X+SxebQXzSomfoSvzYpMba8MitXl9lBb67MGkfX+mMU
lc+xwQtkzoWxOpU9WErCl7i9Gs/3liDaFGJul7iXjp4EGWLItfZFkW00DFDNcDUY
UjGypKEnidEwaPjAS5uNRawiKT9wE9xmo81AJFyj2+PfIMkgYnw43xXi8sK0q4WU
p2exDd0c89WRQmLYZv0aW9k6CR+M+TX9yOhnGnDqCcf3XwoJe+RwPJv7G6KaCMmW
klPgmFZZfRln+yrso/Sco1QHyaBKvOKinXVnrBKMlff3DlcYAA2TzGjAvUhCN53J
KaxxlNXd8SiIGQlstMm/Apxih6+dzbAG2gn4ufNoiRMrcuXckNroyDkz0ZEJUBdj
k+uUNCREcJ6+7tB7ZHeKBBUYeXWvpuI+JIOpC6znKjkG9M9IOwHcoyQjvY7TFJOV
AEgKS4CO/2onSrYTM6bQ6bfkbJTxN3urTjbcW8O6TEnQpaDr83OeS5KRwKOerGlU
ma7PDMnhpVfIhuSqk5kMrpQAJB8Du7pMttDl25dv38KvY0eDu42EZozgkXhAVlu9
8xWR0L1mY33Dcxp60bWfPpp9nDfYvrvI1JMdM1OLh3SdFFfnFtQFFihfTQuSM4WY
uZWvh5unKfbvx34WiRLaAPagEIHMKdfSR/4h8jOvOaebgbTzu1M31Dv9qvbcFrIA
X1P9YeRU8vmmdrkbC6o7xG4EOHv4FwxZhcDzP8P4Uz6kEwSvD7TA/3U+LfBhdFQV
E+KZcpY6qayj6YjyeTU8uQzAoXJB6dX1iksNZUc/7zEcjZWULk34ATj0X3zDFBVD
I6hWHDzJBim1newE43jeYV76CaNxtx5pfv7Xw6TPkjGYfj9pF1tyE+5cWy1SllA7
dGP59k1y9Vb1u9sds81zIaod5QYysmBXWGn3P/pElk5DnaF8jIUyAtwZFpK7Nrjj
o7OqUxrui4QI5mPCOYZmIfeIb8MCFyyxEQvfFfJR1a9nHYcBR6JhYSvaWd4A3CSq
UPc0NyCxkUi5gfcZSHFHReXY4bC6TU0DNxIAUgzzsaKfkrYHDLyyITkqM+iymdWf
X6XLrOQhfWYJ8hodlE4puknYWduum40Pr+Qz5S5+xOy4xyTzIrx7eITX9NwKSOM+
t2V7xJPHztoGJECZ7EAd1GmPZrGcIPK7OLxvm1c5hafPPvoEsCubjkh7Mb9Twwxf
crbS3wu/rLhWAenn5JGo/pwCHJIvwIuViLYvp7enOv0mcJ8kEVU7fiSSrlZpagJH
4O/nQIV//FdEhE08ufasrwPvTOgKKoa3nTtVpAKEopoRzYt2xHyK0kRbbPe2Z+A3
h2HL+vyqWmz8o3ZUyZ3x1H9tBHbLuulQYV8Eq8acLu1ebLRHgR1doDruTw0L5E78
4nyQkbT1XY6rleOv3vHi+0ocU9aqecFrNXk7vlgXhUukXV239xXTc4vAcjQ482lB
RVDtElYfMzwRs5WoMByhIVhP/y2t6FZ7tLTcyvhSNlczVgwLNYwk+gfs28XsN6n6
rnlxgoL8C+uzKw0K1NP3OpSHdJCeZ31LGgEWckXZGicszjo1WY62Ygj9XEjnKQP9
/tqb3jXwwz5OPxQeGNQRlKWijBzmwLO7ytwmXy/FNo6ryTfd+Qu9LhkyVufN2i7a
/B/SyIa8l8dTm6zVRHkC2niyiL+Ur5MgsFZe8nR4mNqHpHs2R+Xx6pxDUfQ74lbT
mrP+Emz3bzGNsasjiwgbj/AU0eOsDKHh9X/3zMYRYQJ5mns3o/piXO7TQZqsskkH
FWen6hKisalYbr+Js7kQgGIovH7ou6QjhsBGpiiKx0seiX/+Oop7m1m3SIEsTC9W
VhJXvni77j4XPFQCNuzngFaYIgj3gEC+fgxW8/9yowvpDYgk4xW500M+vTsX8WYj
IlVFqKOB+8GU8emmabfn+rHvk0vunEotENP6icNy4z2S4r7oWkacqxwInkrGKyh8
Dg72oTjjzHr6Sd6gdhKDoiKay1rHU3yfulo9CPKNvih58INhHXvoNUC6OnxHUxsx
i341RdoOOzeOmp7Mt7Lp+bFJ2WC9HjJj8bkWoEDYtXAOIJQEFS2UkbHIl79+OfcJ
nfsEnzpgNqlk0hcoYlorOntabjcMpzc00SGJhXd1AkovazEBdglm1dh43revTEXa
bMD6R94bTANobX0QW+qS3H6+CHY7utwWGyziEzjTxL+7Ccd4Xdck+kWSdBdQYBVE
Zudqa2QVRPjFo+BQojJnhINZeDM1x4GKM0ysYLkua3wIdB2n255r3pay3vV4ohRS
MfoKyj0jty2VbpxBYnOU0o1UFD1IQ3mPzl1+TC3BptLc+TL2kDyap0UKs/xzypkK
duPwLDiE8nEKcDC54ox9kfJPhZ8ZNVo4w4rkZBUNapEzc1BSu14GaUY2ZtpvfesR
0dOKp8CDXnH3OkhW3CupTfEyzhrbcRXiFHgIpSVX21KVrAX4dfC1z+Pr1lHmVKDW
vKEhDQRNg6xxsdIGKRaK7H/mQsD4DZ/tvZ1IVd376S0FbAP5MA2CA/ml3s+r1sWG
muKLFEFtDSB9+MB5GtMt4PQmcNz0LKBBPXHbt+/DEuKuo036pKik6NAh0ROG2/1R
cLETW2GChLlxRr99GAQdMmdPBmZf1ytwCnML6rCM/WpGzVOhlrthG21gHpvk2KME
MqW0K3wSzOGOnDMGbWxDa1RX5paL1hlamytc7V2yoYXp2Qmu3JXIzXv+ns2wf32b
eKLtwTyvdpdfG3GHTD0h0ZG9z8rzx2I/n6YaAdhYuormZG9Ioi9fu3ZA252PKCNW
ph37FSWh81yVQxeRC1NVKt2cXbO5iM2LvDs1nHGXddis3unY7QEvVJlnGHYXrHEd
vDH3HUl9uN9DlxlLlkjWtzswwNb1tcNnrc4p58Th7wLo1iT1BeMXVLBFjlwWADtA
slZNcdbMBRZXiNAGX/y2ylfWTNIvJ0KJflktRXi9Al4RHAj9ea0F8E6oU+dzVYfi
/M1ED8MfbXrpKXYXHb8gWEAnK9znmwV/AwZ1o33kcHEq0zLXTD3R93OPQqKk3Cp7
YoIDmY0sK+b2aDSnrMZaK+lnK37aIWM5W7ACgOcYlf2iTICc8p9ntEAqo155N+A0
L1qnooLGqe7deC7KlwJ/JxZbaLKT+SD+cW9R2AjfGKvcCFXktNOi8lAXRTWOeMdB
VBnTpQe5hRbix35oM996blgwQ/3C0EAQFdHh+hszDbrziEVymH1R01YPRd2Wgl47
zNuakrxF4FLarceXWA0ncx7SHn44Ov/2zEd0/feVRRCBSgPDrlz9B7zWm603s0Ic
fYHm8odScQ2HDPDNRluWrX7UB0yqPC1k/Lq8BQvdAU/9JM4Wl7guiTOW1715xQZL
PFRpgSwTU7K9jUqBLoBBzjr/IFA/ostKiubvzEhkuo0vmzdh0We2rNclyAC4dbfS
QeNNU/QT/PZ8wpQZ5Y+ccuTOf3yGDhpXMZVmNpS4ukTxzcz8wWXB/k/581JhaOc6
PNyWY6E2qsUkMxYP85nBvQUsrhKADFk2kGSmOykGza1LxrOtHCVP0STuucHbKV7t
ENbo6ABohKHmTBHYjpWZmAkaEGT8otB4ZGAuB0WhZ1WJDgGnJl/Kdv/yDRKGLVB5
aW6jTnkaSxOceB4WHA7sasl9VNtDRDuNWqAmKwvbyNJrjovpD56HiHJCIzVVtDXZ
2iUJF8vPwThEwiARSJZtpZokrZH9JXBgxFu5v1slfuIIR5ouqxEM0G2GdapTiWMx
Euosh1pM9MpmS1W+lC48V7MBXkJe6CNEfLUJ2mjBLPORaFbgtoO+JZuETkLNg5ey
XxUghZBkbOLaPONDh3gpaLqnp/vdH7BShbiKkIh6Emsl+5wg9m67a9q4RO/vYGjv
fehaNXF1Qvc7zM2xeFwo5v88AZaWg/eDNL1reNX0X8g8duMUg044/1bba+EpdHLE
KGZVZ1BDRxWPRP7GkIXpnahfVy7ymW5Ihi0TFuAXYppf7af/oIh9e1+y8yOfx4ei
srUZhhNQ9BD2FbFmVwEaHVAVqESP+82sB0wVO6JzX0DHDGfbDVPQhtCIkM3fQEiG
Z8+jOoRZAFISiT7GSCKjodYT3KmfzdoDhMeUc86GY0mxGLatfsy0wTuqYSxQw4DP
b6OvezLIo0O2J+WQaalup3gMmYGN3mQhxIRLgsCCwFIIddM6W9fBGoTO1adPXvkh
lELO3Wh6XR8P9eqF3lFcddOoRpxxA5ZmtdH/TL2Noy6mj5Ackudg2JqlhrC7DkgY
UY6Aa/S496meSvNp5uKrd419ijy2Z9MRo7y16lMbqIWeiH0v+1SUmuRDB1fWUbB8
9OflRM4JItQH5SaYSdVetWtw+co+BHmbQh2rno7koFO/XgcgAFulhXfe3l3o8bLy
IQ+ZSGzCXZoadt+zzowLOIBK8ODBxm2UR9E7pjKjfJk20tSY1LDs8T5TDSJEY5om
cFHoIBg45He2fGk/1sVWvmTu3aIVDD003QWkubogRauC3DCVvgbaFJac0ZwWBOcr
fNJZTLc+Tsf56gZ3EgRYf/p8VN877SoCyrWp7CEiTIGQDsw5tt5PgTYgxSE+a7ZR
xZthAzR6/gD61/IhUmZirFmeeNG3UdsIXVG2y/imVminLt90uflrZlyHsQw6CWG6
Nh6MORrUHW9ClC/1OnfubALVfaRV9Ok8E0cg2SMaFWCXz22zPZEfOJqnZlscAbEc
tr1E/XjZASyEBatKDc57kUpXtoLVyZGXRDtnKL0HD+Wt5IRZqB8ecEa7JqFrgbP+
5qoz62gN1R4R1jbTFyWWz5untalgymZrW9z7u7ComWz4ZJTBs3nkTR0jAj8/rXM4
GlkQIZz+diE+tqPlO9e5Dx36dXHiTeN0DdiQtMbiXsmIZjvkiy/dmEY69xBc4gaL
bFprx4lP21h5JqZ2o63Y/hso9vMt+6tH3ANFG1KuchzrFWAAvHaqAT47meLdDNLU
/zcmQF0MXb2Q8/3bV6H6yhYhbbzR3EVKsbGBWrzkSxlN1vKWk7Y5OAuKEbh4Ir7/
3g47BwHwLE3eT/OECsmse+ozrbFU+cG7p8tQOEse9ggb5Es7XaYvu/gOruJUT67x
uiZ6J1wJUtucAwg1Tie3hv9cAFHTcGHTjelwqwH+bB8wlV3R4u4ETSaGwGKGtev0
p98YnWWebHZqFAlehA1KV0ZHcJNMHQRvHvMzd9BXWb8HJrWMVYw7bk9qufdYjpnr
l5WDZlC0CyZ4lv89vLiJKFZVcwer06eRpgMSlzheXNu28LWhmRY5tpn7zxiPCSK3
38Dw5a9zdHW0N6Pr7XcwQT7wR7x82YFsCdfvlJo1Zn0ZvMNkrOxJGt3v0rwLV2Ol
3vKOueeUhZJJaXtbfcPtEtu1vuHb+0PDcenkOUGhpAOGP9tLZwTkQG5gm3fluvNb
Q18IMmeaShJoBg8P9p5Grz+yqTyBdQf1sQkz5tyDN2rJxJaS3rpf8ekJTxWkvLdh
EDNH//C8GkjS0tXYLzZvCK6ZGdz7VZrXzAIHUO8igU2LiftYg9FNAQXmEBBtz1kD
hJ9sgDay0Np/8aVpfaSh0XHnZ13ORySuqFMSm4CKBxlMUt4jQNR+AVY7B4euv4fl
TIoctnTtahJWgI9fSW7nnlV0MMi+3UlULwGishbnNFFoYQOYdP2J/ExnQBKpNyDp
b+Z+XvJaZ/FdkzPgbONpPvLYCxiD2JuznBa/DI9uMNRfHSsWvOR+QEN1l5o8khZV
koJMBLYfWn2pY+7jLwW1CZvxfono3RPwj0xEVJoknFgQOcVsvTXbnKNDx9jZG/ID
81jAL/P6rdnvVO0r/AkKSYyOfhzomvR/dKrvaBXJF2+uiuI8VReUWGfim94eGBCw
S09+9bcPqj4uA7FJYyG/o1oxJ0HlrnMcQU0VdovpqV/FtvutmcUVFUih5nhdDQrd
w77/0nnZQGe1bJDCOj3+NLJI35yPi6qNYjrDZMyi7ceDJw47Sc6uhk/q9wm+sQ7q
NkTObV9LUY/+fLr1yH8sn4yYVB+PxhEUElohq0pcBPJquI3DRBytU9W0KpMwDO9H
e8AsOP4rdwv1YFvwkbWyDalRvypC52rukSpW44HcK760CoxCGlpwefOp1CK0oy16
UPGA9FeFrTmg4q6Tg8XPvbwCbpwYNf8Qlw7hkwixMpgoRnFashoMebsRrftbEb2m
MnpIGDTsnN1zrO2s9YG/q3SmjR4RF5HQSZdtL0Y/ni8OYAb5sVUYVTCiQ7k4mWoo
smjSzKb4G0aSVOH6hVUpoqgza1knvNzlR/6BSTzP/T/CL/jlleGbxO3K7dWh0MFI
B98E6B9DgxR0NcD0KDfIDQHz1QUt8atVs885fU3wwOqF0Vi1UHgJR8xWudAduN3/
ZoirTFz01DhYqHPGsJ2FU0PTDftPNauRA4juGkW3ye59OOG/MSluJ0+F1WXipSAW
LF56geJSKrFmvlgyr9yZs1YZWzYqtB9QYZ4r60AAtux2Szw0Ixdwl62KJUywVxQu
BnOYIfELyvhHaxJ9fydzgT2xaQoE7FVyKk6Z69oOeErwTZ0PrOj85+Wu0VOeBKBt
ZDDyRPMSwFc+Ri5dVM59ACMqjr2UwQQcJakrwrvqiP5lJKYH2KY4v55NqLx6fgRM
WscTaAFo21ATJtJ1WLOagqEVxTE3G8Ft+KwGoUuC8XB8cTXSyTosqcLTtVv5dBED
XCy548Uro/KZp/PCHcMlWPshGdwLUfLnQRyJ0Pbt1e/sD8VlOZzxmvb8u4ZfLL5X
nonGPFluk27xu+EBKMCK37IX49ni0e8JgpT0uQzrpd9z1s/3ZBQdezWZLApygHBI
hW1pR6DlepheoVTATqk/GlU1p+73p9D2t+USRyt//rjJvS0NXfiolFsjfy4Pou2T
xC8KEzWX29UWk7xxf44ev7IsvJDFK7pdZQkdmoWAW2AMEtE2STcH6hq1+0KnVslp
WBrttAaNMSfuOgbTRSRFVJ09itCjbQorVJiuId2BVZRxrHUUf36et7QFQFs0IjBZ
mIoz5iyyBUetcNH+DUbxpfUJwkVfXiGhKcyuy3g56lGLnuOMX2tkZxYJIW0nAukG
SwgPSereR6pclk6k5MQxcaySUhRQMsxzXu00IveF/g24w5wWeCmjFHStZ9umtOeT
lRngF0fM8s3bSxp+2Kwjiei1N8Uz0WU3O9LFy8TME0NNPkr3zZDJAQ+DOusOltCJ
P4B289oxCvMJ+tP0+xOYWgn8o1nGtCIVPw9h9JdxWzP+cpOtPZreXupoCIg3zVoq
Be9+kLOkHcmBXPTK4XUI91ng66AdtTrv7vEjevNV6ufHjnO/3CdH66jswExhEQt5
nEZmhVwNy3zTwNCU6wbfDPZbx7z5VEJSHq8d86E0FV2bkztcwFu08KfJhcBOcHvP
9um2d44GTFL9RmUG94qN7mJJfkInyUGsUbijiIuicvCdX2AteEpKdne7y5QCojsx
XP6p9Knh6p8aKDmi86dMwlCIkpaffzsDpoGXlSUiFLziPGdBut7TggHJwEsnXwyT
uqpOiRCWEZxFQXTaMqIHq8Y1V8vQilClCpLblguoeG1ZXuVRX0dKKoInrkjNJ8u2
LL32tCTjAoUGvSs4rXyoO1x8zOP4rkgHQhj5Y1Mr3rtt8YuVOSUwHbZgVWTSrVE5
Mm4oM6kBK879STeKSlgBSxHBHCqvDMAdXLNWmpMoJrVQl/kn1y8y91pleSJ18dif
9dz3riAq2wkR3KVarFINIoE/7y9HQqXA/xtxx4a4K+V77nS7Y1Yp1bI3uO7QlBVg
t8Rcnea9pF/jydeRadIVASXzZuRBb2zNFL0MLeTv+hw=
`pragma protect end_protected
