// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:36 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Wy87d62aWs+iT0XAFCVwee75Sha2d8yvaZZ9/O1+seIMDCbRspayQ5gRHsUt6Bgc
bfJEABdC3ckZxJdYtBq0Unemmfqq8uSEObSM3r7aE02R4d1IWWPDw6IP0CSnpIey
V+JdSVgRVuKSc9eP/YCe1LcW+xt0AYYJOA61uuBnlwc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30848)
MsrqrZyw35rfdri0+WLw5JZ3hCLafVtTQL8PyKypNjYMUaA5auQJMEx/h8mzVY3o
7tLfwx8/YI15SUhll9ACQNTV3qLQR2KHgLhsH0xqMxMkedAPKZPwqeIux+a8GYN8
s2pYjoDyf+lfu0GxBv2W+uYHKo1H/JRjgITgCRaVwOgXdtVN+zbhgd1iQHrQdq9C
ny5C7LONZMwokhaUzY/jJf67WudlkccApPUBrnPllseGcjkdH1DgoyYj6AxTrOQ/
H+pOhlyWODB+d/uhLMuCUVYnJbOxUNTWqLMsVkLKvHS8WiYI1/n2KjvnyFOj62f9
j1Mqlz7dEw2impAz8oVwDLALXVAfm9enPFJON87sXMpxYUTOA6YxzbSaX2QcbI6u
3Wgqo+jWXtCwEmcP7AczGO0+w14p2K5xRVWvx8ZOrbXVMimZF4xPxLgKoVRxV1s1
XH+gqoGGHQYhDR1V2fO6rCwRIw4Q/OR5q0RKDg7c74wKbHm4E2xfGqWFVXkcEMEi
dvMmuCRv1QCOZDnqAnCX+8HZqgtn0bN4w2GA5XA2iQZxU9yGPIg+HQ15W+4IyMZK
Pz4g+XkITwKSoyP6cd148D4WNBViFfBx+PuHkN0DVAITH8W3gUbhdglTq8cbLZhI
rG85Ye8875r5c3M0+uUm5oWMjSxkAgAeteR8P/UW+h/dzDlMQfj0CP+5CN/kymVJ
gbVZm0qbmJhroM2jJHkhw0RJnU5XRdK79RnFs40hUbdpTsxRaEPX+iXWPZRV4R21
tb+cpI0hUv4+FLIlqTRjnbnFg4R4WEClY+0hU9U4PXL4FURkr++NExvsCfftzgtJ
ac2XUCcIsPrk8zMs6/LG3NesAatV4bcchYCkuljpgq2nYGSvo0tss4xUISnI+2u3
BNLfEPAHInbisiDexG6Ga8rM7hGAaznTd92WGRMWbp70YWRYPXjl8BgjMkv3R2OQ
X8lE6Z5l59mgKbUypFabhzAuF3kARC1LF1UB8Kru2lgltIYfbvAsOKuswx3m0ShS
iaEVg/F8FgvSQy7EJe7TqAn7zvu7oWuPkTpi13n3rWtDsHAXqqDJ2cnWCqTUWozQ
/SVKDbmrAQDiCnlzuhsb8WcGhpKrto3yLrXHVVsrQTxwccJWX9JwyLIz17aaHM78
kU+Kf9x7sZigibvBAAh038zAjC2JT3UA6lKhsAc+7n+jT/ksxggrZVxYIuDS7bxI
axAERKdOYgTT2+IhYXJq3Ryl0ClVI1/qneld4k2THI0Yp8xJuNqMlugDhYsQUSKh
2HcIGZehgQ/u0FihAxSZ8v6dnSyqWk7ScYGbEtcg4NHFDfM0Fa4Cx2rpSXAh/aGa
Ov4cisCSvAkF0NNRPErlpWYEYx3kGoSGGT9GpWGEQfy7E1AyO2d50zlsagHbd4FP
XD1MakfjRDWZd1ZlituDndAnnoxO/6bH6MkwL8SR1WXhHglJhf53FvFT9WSCuEkM
JV2RPec7fiNQHV4NzxPqP3VTAWMQ85HXNH/uyPFqhKkwnFZSjRCTSJXwJGdlSpXT
lM7ABKzcJTmuzzUU6JvGZ6fsS20dL4p4004XZ+pLP/OFQ2Ibzj3b2jXfkHwnAAcN
u39Rzc2RPpNaYqsvhJ9sRCH21/Hrrb8esiBwfouBydH0h1IkjzSMa6DwkiI9Gok1
WW7JserkCneNpwEvnQJha62hVBJMTLfBCY2tD/l55nZUwhxzcnkuj59AYfebzbam
iz3vGLbkzJvsJJYT1n40VpEbS6/Uq0tyVwtz+4DrWUq+PDCHbBHd1MiH7PaucQ7i
j4UT4IQo5K4sqzs3+sKxxiBitkbccrFICokBfJ+1JqIz6nM1S0SsTrVuDjvRetiJ
mfeIE2aC/dcRbR9juLvokVqpcbT7yHZpC/L4m72hhhqKknVwDN/xOUm9xWegfcVj
3sMJYoOCoHuQ3JQuwxdbSJ3HLoD96p25c/ds2iBjALHIVvNR79KRTvMTTr/78Y/e
SyF8mLSdX7kzcugyZ4+0dNZ/bNOGYbpmARs39rpfS8Uh/Ffu3IEjfMWSugrw36hs
FD8zuHJPHaX40EmrzOds6UlyD3o3rZzE8L82Wxxaozx7ueX84Z2Ri+TQFUqlWsV3
y0pARMbqJMI8zFLP7WiWSnpRi/Jj2c6+uGOwkoac6K2xzLOC0xiGnEFfe7F/jd2y
gVxlhqCi2y2OprGzTKCUwiqgJSs628igLY3Vg12lSGXZAF3uq4GtrDC3OybApXTP
U+meu4U3MYWQBZybTMEiX59La4CIYPgV3bPppupWDr85sI6ccTlWVy4jMxZGjJiH
d/t0PN5DUDIefewfF9Zx5pSkGPNLoZT16rW6VPpN6bk6/31pDL0sK6hpx0c0oL/z
ddrRsmo8plOc7Ntv6CW5AjAtqdmJInSTvLnI4DgvFNEOzp+6QUQTV1VCr4q4ofQ/
Kc5VWBfvNMaUOv5fqOKv9MmZdmfwQsFauJQCOz9Gn2JRGR7wUhTmsUN7toIzs+pM
Bp4gxxfcZtBuPrBmKMUV6mIBUHahoXW12osFrJ4wHGG3yggZQB/iytJXht+r3LD5
FpajJMbe2L7u9SxJh58wWlCxuHMsKAkN+DbullAg2M12Z/lRXHMg1mCSNWbOVtzM
n+0ntBH8mM4Qu4CefjyA0E38dWHUsYBTm+tFYbr2YiqyyfU3TvzFBWzs1X6meN6K
+Fe7NsNVxmvgspGjWZuGCY3A1PNgbLxcW8QI822tABziUJmpvki1i1hPoBvMN0SN
MjCS3RVQJECHKcG2y9jefoLNgQnXGW2FTqtlAsQlIJ34fwBo9KcHAmafVq2DYT9g
l+Xhh2nTEZaQ21OjgFNc0EXYI2NCB0Vcbmm5rQXRlqFZyOZsZFGahpc1yKtAsKcY
WMYQ48DCagO2PlsEiq0+kyqha1cvjG/iVNC/FpD6pqsNm3Z766NJ3FSTkZN5qIOO
VzNHjL/IMXpW/4ZFjUf0khTBrR48L3OXmJOJ3jPy2e+2njWawhNk3sxrs/LmtaDL
f9x8LG0bS7pNFtuXghQPrdHPwaVzxOJmGJkO93Rhgzb2i158jC0aAXtiY2Vg3gjW
QsaEBPkgWVRRTdXRygKpzIqPcyx7gtsEjVBPB3DUzukJJWIs/nOcWKcNyaBgCwP/
JmDxOf2707If/PPibffi9ZPN327VN6HhuD2nMNOWtv/aUMFj+qyZbuEDbFW4KWEW
LLkVoOxQ9+VBuqn1tfeGQf2oouw7U2kw11UbWRA/ytp4vYTjrVbodFFmXcg3bMBF
GWVzSzyrh/lLsb/3dZiqqBNUYeqBkpr/K2O75v16ZV6xB6hLMtWkd33nyxfoOvmy
2g0z9p+sezXNwHUYlIYjJZpLJi4LXsv94hdNbcmD6FR/80Hev/9sjXEz71YUO1Es
LxY/yko90eHyHWXGPOfavr+ea9sjApo6D1DdO86N2iny20WzNUk62K8G+C4s30ev
PTBmV05OpKo3zf8UtlttN33SPmM02pmNq2gGEKSZevHj1AZGFPvZlA4pMwZ7lBpc
MCxCEO755qcrnorNLAzI869MDdljVvuntp3KMWLYffDcnuggMQ0VOjk9W89gPfGH
mqmErME+AUh4VvMHTSq1M/u4IGL2sh4lMUp+tm4tDjBwIFZC1LK/NhAFDr+MNgP2
wtD08LWux4Q+kVjlLIIlnRggTwS6GPan3QyxKdJo+uL5L+JElpu0L7QZis2WBzAt
qyxuiIJd9xVif3W2SqZFIEzmTvnLtSMvFY+evBYlsCTStElOjaY0n9AoxzuF18tZ
/vw++exEnyIr9WtN/qfASXDLWG83fjMVElJkXArMjm/UxTHnlDZK9hkaFsKDJoWa
Ljc9RAA5kCDO5uFtesQ1ciDa2IdjSazrJygbybzFbg3/Ewpp4nCL8FO78mNJ0wFu
RHHlvIbpmyuXXO3bqvukutoB7NvO6LLodzOrmF5822TBF+TOdcI4BQFA8NMGoWlM
k5MwuSAtLuQa4WyGRHQNgaffinqD2XR3lJpgKZJaCPPsY4acLx899YZd9p4AUOA4
J38oFuo0v4OyxpjxIiU2B62E9NkIyHKpmaAwrbwLa8lOq6iRLUzK2tvevESqnv2t
RArr7ZcEYLB2RxROS7wKK3Ro09OkWAe0fAdqgV7VUQ4QNUQPA3Y415NtaEB3bRas
7dyhQ+2SWbQXSfIXswCVD7PmyeyqtaaXwqdrfi4eS0blU4jaViysgEuAVssPC/r2
k0dIyEUE7MctDICQl96ELKku0tEpdX8MBOMchGahcdTVfnT48gLw4aGEXCuyoH6m
sCTNbhxAwM1S2HYyELsijqTlhwFczQhYKQq5lfTAR47gtyYMxzb2vPbduzmkVMsQ
4miarl3crP5yQT+PdNtRdOA1l/WC5ByR3qO7PQXDyKi2o0rhPI3WBvFD5YFaXRNI
FBysocreexAd/1RVNqCxM/C0i8EGJrla0EkQzoBtLaKM5uNBrVpd85JzqKOTjlJT
mMxAPPeA9vDLnK3/bK1NZMYjUl3LRYCmWKBPrRwDOEb1j/8uEvvqUEqDy+jNj8mE
TXxyEiA+y64gaoFUH3cCzevKXWVA6NRwnki71q69OMoJjOJvf5p65fQIpz8UtA4b
YhISYIpach71bYIUKJlV/plnESdF5p5ba2ugPGnmq/WmDtmDek+CQl+2FUg9JLVE
h3X/3ZKcux4YN3fZdnIpi/hCQzDLpSepzBG0g4sDFZbgp5FORf54E2kgMJrRT1uF
2fVwYnWXO5CoJNFumVnKdo9X8/dUYAc/jCkIxJvtf5q29WVXHK/lKIi1nGj4m/of
+PP6jQQyajMBCsS6z8/xTkJ4OqTVw0zhNyBajVSZXBlNkKOclRvgMywFMpMy58HW
WA+kHwlDqbQmEPUDggfCn/tgGnMgsTsK45wdPk216+pdotOGuF+Mdno+kdVwQ0FM
F0/yng9HmIuvSJ9FzA6ZeacYhmRT7NecBDCqLSQq2kDrl7FN59mEG2kMkDMDT6Vg
u7njaoF3sCF7szSbru4biJayvvW8iTaXVURnBjlbcMstsu0BgtKB/xjT6CO5bpEh
cZ1wSm+gndu38Ni5ByQ1b+HQuE6txTzqNrOmnGggoCSY9DvQFTTreC9a9/lmuImv
j2Y6MqLdBLdGNuAd3x8fHzT/PvwEpvHvMod7izTPtn9Z9JI7KjuZtU0733uu0m/4
th/gkF+mof2V0d6OEv2DMToOjDCu1MpET3Plt7KdvCQFgCnAFtP/ycA7MlfIXdaM
b6DRrL+7faJBKc08Y16BI0q8JCnV46DL7iTbwylohUenTumqwf/qhx/M5j2xUgeC
1DZJBte6tmeUWLCqh9+xvh5agJSY3Ae3f8wOCieu0jht2TsNZ3GLbkOpbojQzgLS
N4ov3LPJjLaAE8xle1IVGth5w6d80SVBQAgUC2qYqFgzy//W22GoBNYGHEeF+2lP
jguCCYVIHdG7SuwL5sxkYl0cNpdX8R4jMq/XfSNgrXWU2DYGDKZZyb7CDl5lJnv3
UPGQO5gcs4pj+c/pJKWC4TGDiVkhFrbxvEPwbJee86m8Pm3pyPHSDGeWyYBbLwGq
lRXcBjvr8pqtVHxI67JfJKvzvYvC+cOg0L802nIfVkVyRl6gbTzQSjGfdvQl5QtH
R8TlJWjd5DrCnDCx7Zn6rwspEyDVmdkFqTlENajyZFOFYit+svTD0j3afO7GbG5a
0X35oeKEyF9KfguJVbTZ8GQ+6GQpo0XMdwfjtwEtPd90OFgGhfC3FMwPZC4+BfYb
8mWxA+muQzNCrCWNwE66Nxz7PQdGs5/JHiz9m9KWRym7u577fEN4O0ntE4pUaXwv
MvEhOQQUO+WXexGJBVrC6Zd5psLByJrlF3GEJGRFlHpOdg5XPIgxCrmg2wBhsg6U
TqaLaAR1UUGCGRzkzrvimOy8EzmmjWunYxZ2oTUwZEerDeQZYqL0zbmS7zIOzplC
QVppuktOMXfU+JGgwtGYJ5OXwJ5zExwZV4ADPrOPoGx1fm+VADlso3J+99k4Gjpz
F75f8hw69RBhXCz3ENkA4QV9m82mBgTG1U21QQVrvfd/BFa+f7IlDYANf0Ar6Z0Z
OKIhxNeoBGfCk8enOUqbpYME9AIANI6ZyS7nr2/2UCFdb4NNsqLFiU9G1JgcIujO
5M74yNyu9Adfu8FlRUsVFFFs4vJyItl5tWIIz6vh3jTz+ztXNjOw6g5HaWpRELgu
KuKoSahMxUJxqP87ZC73qRPgcGc4qmZ6KHzhYj961z+c2Ns35bwduBgvUQVH1WB+
5nNJtM/ySBMXbjUu8ltE6VHKHJOMKgcQgg9Gr5AziUOOFZP8O5PWIRE2FXB3nGMz
j6r3K48rCWJKQ/EOnPvpngcrznDzaJfxKAuCOtPqb+WzqXAfYgaV7ZgBb+yGc8oa
n0pBtU5FPPmxsHYr8d9CfQlJ6fyiO6DW3pwLAny47YYmYK1I2MoOkXh7Q+EaVFJ8
WQv0HbM9WHltfhelWX+mW9kGiL6KQXgUuL6hNoOWJA6x0Der4WuAlXUZtSFfuzv5
CHnTbt8ekMFKg2x2N9jNPyq15lQfeSdQsGI0sAxrpftTFNeVh9y/wLMVeCRB1elp
rGsBWz2yBgzLw62iDwu9oWfhSsOVYyi0ja6g1XbozDdiW/OJdMBPJmd99AqgniyB
y2yZvsVwHdfPDn6uwDqgpEpdtEL0SbC/c9RBjYbblAP8T2U1nte3rMeZX2LQdYbQ
xjAYUlhFieE+CjQEfC9Y1XLaxKvhBgmXEFdow+7vY1I8y72PONT8d7ARyNviMyLT
2sYhuRlxO6oBkJHTWrvXAtqlxid4f9eLRikaGvTaeRJ961UwL1uCKD0dN4G9gRCj
E2gy200ASOTB5B9yitcYfQL4oUkriG4M4nLVPn0tcQSy3Zj1rIBArVjdmBrPNwCV
N/eBUZpoQPvFh5vkLNRz9ZsDfYhL+CQP+rSP/doYjQENFEeKSTEEJwuxeIF3jL06
P3Xi8xlGida9PcdJR1JzH+uQTO1fyzjM7l8feRUFvhy7Oof9LLfpvHr05MXtD3PX
80nWBr7e0ERiK3HhDhiBfjt0omyxMjZBucXmzwy42EQsCmgmGokiD54xVS/ksOGd
HOiFytO62Zd3YT0gVND6zMrS5aNhlZHCUBw7iomv9PyUShFVgkmAxKWrchSMsUYQ
tcY9nIKUgn8aR7Tm6BmyqpT2S1ldkqGzoK/mYwDxy4KEXQ9P2zjy0g1Fi8JyIV3q
Jq9xGcX51bAc+vAkRbw869LOLCElntyXKexSLSwvs4C62ebesAOyF1yDnuIbDCeJ
++tftXrppvwN5/VIoEt/zk5Yx0NusWvTN9AOBfKHmTjZ0XyODgXtaZhMS7povFUA
wNwUiZcHIWHzN9W/FPMFtsvOpIiNW7c/1865Injyb4DZ21aIVg1hy0cVkCdedOxc
0LuYb7CGaf8q5eZUrmaSA0TNCQmdTNBUHozs33pJeUaqwx1r0sc4l6a7j567WDJX
pS44CuhzNKBpWyLp7PW835zjVUJBmxVzOqYfID+cTbJA1FI9ijCLFodewk3JJ1i1
MjYf7Uh8aE5dy611c5AQ9IHJZFt/RyeFe1KNC11rTRVaLTPWfwNGdvXqdkC578K2
8/iJDgru7dR2Iqk50Dy8KNNrinbx9/hCkAG4Kkxt+SRs8Hpe9wsoO5GabtZJ/aXV
YVF0aKrJUypEW1eO8gGENzrqr9DqayzrpHsyCEKK6E5OLLtzJYKquP4tLmtqi+kY
6v+jcrn3zVGoaxGBt4nRmJpx3IUyifECixxY3QHeLK8hZHLQ1MmpihULDqCrpE0T
T5OWGbP6vOnAb9780kkG/RfunuXkhF7FjOuobBfPEOi37JwEtLi0WMet+CyW3rEh
DnwGfkLiID8Y+0ACWUsnyZJuSJSZdqcfPxYoi7FPH351dM6U1lqLXqRAOS4cpL0Q
Qkc7ACL5lS/yGBjBS1DlaAA3BGMzu3nkxLe5cFDBABDuawPMuh1HvJtPAVt6FpHY
mjS03yXw6Rk97b/DqOPI/kxqC6hznFaUJkrv3MU5zAHJZ8BrHW4Ev2jrUFc0LxFl
lKjb+ez66srZIMW0+DYlx7hpVBvYNaNaRtzHWvA1PzRJQo+AfmG9fEICFpb9olv6
IWDz2wcoONf6RLFGXd3zQAMzTuMpIrrBjadBT/OUhL9aWbFZZ3Ak2cGPGSWq1hGN
y4XsJZzlAjzslvjZV3vzSx5jSmlYKSy4Ba02zyIK5rNyjLiKkeiL0xpYy8/fecU9
bdi12F9dCRAwdb/QS4LnZinf50+kNxa8J3yGiuwSYzpO0jcA6Qp9eNSC8d9kU4Nm
UeoXCJO/fJCprQ/LX31q8XlunYXHmcP4NOAdQnJyDF31/UlwyB+JUzuaClj+DgZ9
+Dmh8bFI+1pfUOrOwYnBqSykQXpKL5nDcBDEhc3EjFgIvsB4TTJCEQz4el6NTo4U
SOipJssn2NqxNOwgMLuU2TLR06V9VFSNkDUL2nfN8C0dxkO5ts6oO1A0tGM0x9Mv
UBsY8Z1Z21fLUk7C8mZlfUaCMU+qT25aTXvxkrSAhuWwcecqzI9+/EMD4/8bzNJ8
3cTCsV2CbKspErFB8x38DseM44MI+1ZaItiwAa94mL7osQD/SzyXuNWKEAF1Gf1d
76Mq6sXA9rHRgBk0C5iy6snjlqUJGLlGghqp0/CxoURkeg890lP/d8HjpUmI/nYB
XoSiYwSdQKXddHcmpeg1T3DDUFdss0wR9Fq254f8PvwvA3icra98BS3/INkXSyVg
InXdry9dLf+XfZRau2Cvsv2O2bOJVyxcnRf8ehJMF7n4X9/+ej1Y2UbR6GqkstSv
xDsOGXdGmJJfwifjP7Nhva/9kB3nifNmAi5wPttXMV+J2GI/t7lgsSu625G6O/9p
SEoqqadpCjjxhSdc4ZdGZFJigbeSWiObTV7ZiWja3cNUpsasBQUhzRmVUU/qvZ/v
HzfMMzV4z400fYdkDUIwhygGRaT4R4WIn0TE2xFb9pwEvgSv4UHRRm5gaB79cUkb
skL+iWfAWueVs3CK4wGYRmVoHEpBs4gcNGU6eESP0fPngb8zmzN1SmM428ju2jAM
vDNyHtp1bicN+AujrssSfjDDGOmRdFU0Y0uzwXTroWC6zcyEgj1gFqphyQjA7wk6
p/JWmX+9cC2DlmeyZOlNPbyqVFCfJYmmJtJiPVz1jxWLfa7ecd0VbK6fVASHkfsG
2iJFppmp3VFMrsFBw0E5S+kiUJREkat7SqZEG7ggNsQmn/rzR9DDWxNTS25AJewl
/DQgk1Ldx7fF97h0oKHKdQB/i2CrzcdsD5bovXGmyRdNsxBo9YCKd7Op/6TwbrGw
p5eifXoNt8RUJO0tuYWI9+bmG4ZLHGB+rywrSYMwV1C0b9Aiqg6AP1VbOF++T2Lt
dhySOCIzhoN8VPsMdECPLFap/XVTN6EgHQhnXaKvPYrJRWEGv42D9qfO4/m78uOB
cMilvu0OCzU/Jt7pwyrX1qnaQM/9Maz0HcJ5YDy0g4m9RYJqSh/07hQN0txfsQXv
NQyghEdGhmkivlsX6S52G3LMNeX2vrcscJIvMShYWBT92/regYvdUk8e9och2b1H
C29wEUTSLhW5U/gcjuqH0ux6fI+Crp22oj0bh49FNqQruoLbVZSXqgxAmQ54pNtN
knLbP5vtYuDBFnlCzFD29yxcywIZmQZO6G+r2Qjk33tcU1kY90tkb/AN7q2plNAc
xxy3Wmlh4C3ECgUJVEb0BDa5hhxi5h/EqKUavLuhAhshUwM+vG1JrUxRhN2DIsnv
yb74+1pT4/bV8Tbxk1Vt5qHHLu4QlckQsGa+Qld/YriDfv7jDEpgKRoVnWYHkIDo
rvUnzO/jx/bI5j1bupfrp4/8gVVXGAncxvf36XLNGVyEPMKp92o5omP0wugRhxB1
tz711h4ibqAzH+vJ474I7oPxrfzsab4JCg1sqUCRNypdLb5bgpbpZ7irub17ypUs
Sway7C6NTb9lMW+BZV71P1KbBK0sgGmNyjJJVzz63q0Fpm/RXJU3caej43qaZUO/
v8TSGjCxLAjnOEVummqOvPJkxCqdj6WyvGgnFwlk3sMatLj7CuJXH+hr2MqrO13W
Iq/BFWZko80+CVaBHmZ+XXbOGVRiS94krTNsQ38S5XqOIZqpaYEr7RqjvlBxbViu
dz/k3K1y8546sEDJYh148XnCupFL8haaI6t8VuxaXXGuVi4YagP4zMfQnKtC6JzA
sbECGUv4YBDRC+uL0zq1z1N1essWfIEaR5YKwVY27zou/a38U/UcVGU2kN4sQLqL
fo/8qTWfndBw1XsgE6tfGLdDCoJ6wDSP8eTbOVG2wlnJNzcJwZ6I1vzW/JzdUIiC
3Sxzd0afqrzPLayrLtVK/ujdDRIdkmw0H3iRajHeQJKVVdtU59ceZ+TdGX7OVwH9
vvqScVyzcRgmwxs+fTqeWFlvd6g6h4jZaWnzmyoOQCFUM/mTIswMmbmWSxcOFDMM
iJOnn1x7NgSPOUMTvTm+D/sZ0dL10axRlN9G5JHggaeMhj+o2OO93fPy3Vks7xvd
adMjlPKxEuXfOJQEjf5apQOyo75kf8VoR/jlw+SPRTyJlqycLz8d1uqVQMZp+31y
OM7dLAcI8yD5uNEX5wwd/A1OGmlbypYGit5kZ+aWaywsdFoFZ+w8EYWKQ6gXQx46
UM4KoeOQ7V+AghwaTvC0eJNk/cBDU7fVWVl37CPI8mMwLb44YzxQtP6Hb1akeuok
/7GZxYYx7dn62c0qzQzPfqTK59Ef6ZSSobhFMU4vVxmMgCd3EuAG3nrBKY1Ab60c
g7lHpp/4hZNiSg+Av9W+J7IzFHA+K2Y3XaG3+8H9tIEk3sOZZVHCsC0F9eRldb4V
l45f/kPazsoX+MXjL9WfTqhxFqvn6Zz9Y/HZtUpB3+ACGEu876ZStYBVGVxz7wNQ
g2a3RihmVPrgz/ojT56ZcdYpRjlISnmzzHMttqFCD2GweG7nBAHg8wb9t2yeYnU4
ubqDjvh2BwMbXxsR/W1G+HWgHuLQnoamzssp1p+pNCI5etFq7Us9G9hIT4Ku7cqQ
W1rg6DxwEUdV+HadUVkPtvXUUQcgQcx8pqWJNr71nzIW2WR/+uUgff7LEgxZGLPS
xRF6X6UK7mwUp4es4kkAfQ08WpZgH/n21JzDd06tbBaPhcuKUj36HJvv1K1RYKIQ
YpmTClEhBFimW090df1+hWnwshAVPbmfXqsxNFy7aGAb4Af/WzFnvvaMEFyeh+ck
EfWfLfTVlJk7M/2Sfay4Qd7XVnFJ5zqFmFiBNl3RUtmHBjBazNaP9gySDwv2kTgN
WgbMyCtMw0dpw86/+re6yOn+Io9nwsWeohxOmtHpXRr744fhJkiycbbaEMJ7xmdD
KigvtoeKVduGVeUZ6XgrymQfDX2q1nBnvFGOq3C8bSe7pgusaEsw/wvvOFhxwqcp
wmwrsJgIPEFIBdWPvB/uEc1Bqg1x76rdkhcLZYmsYei/AmbuzmwnOwgBqPKQcP9B
zQ5OqITXA1C+rjgCleB2gMiNC2W34O8LDOdnpKxe8O/CYaOt8L1e8gBQ56hpNqVw
AnIulAUZmDPZpFNHcNcv5rCQYO6DSfjb4H25e4NbKwflU9dAAleY2cdL5ZgpNygp
6uTEFJmYXiBPX1lWC+pexGD/yjPhEESp5UI0tC07/Z8X/H94sgXvbd/by9bapkSi
GLkIrF0Kz6lqHbKUlvd0J7DMM5tlEbMa84pcoTZE7cFoCcpbIzL+S0kOKO/AvVz9
fkLXzJoJSkPxBOKJGE7/hvh9yliXi4/G4KBSX1Xku/frfGVLDCD2wqAJcZlu11+u
6eLNOqZAO0pqJfnzmxtYJXv5URicVeC8LVkZoHpqh3FWElbclueuegf6lF5EFOZy
9b9AEpzA2rb7+nbXiL7O1MnlU1tfkA19Z591XJgHPAtE9U09Tg2kl+Z/KJiI5khz
K/8FxWu/NJ3Ax95S9r1CX5RYIj7/sU+M5tcNNxBV4p1qCGvwTvx8tbYk9xUKDpsq
/5MNRKvBtMGTwwHY0NVVVbvb5SIxnGKn6bdTXQAmsdWOyyFmy+fldReJaJT/ZA6K
fBL56KCMq9zZ+Ol3pEKpyzKn0JAFdRqyVNmPsTCbK5mWZwLwXQdyXGHWV/WDFaJ6
1U0LLP+jsOnlzUMbPB7nCPd/cG+aqRPM2f+keTKnzxjPev88s9za7HP0i/zkK53e
dGFU61EM3nKLEyYE6fJnLQ7NvtGtxNbVH0rnUuuwW83ItubjwZLGN6akN1zIXmPA
HKFgfVLjSjSdox/OMXYiBaHYA9YQmWvybiL6hbadVMLnFtb7JmKrXJzG2FM3IyF3
/ZiRAAeBgaxJFfn+Nf6/sQf9E6SJBx4RZRZ5VCGyIzMOhizLKmuRc+9tKPgetEgN
jFX6O9kPCfqdOxuTnJqf6GXvR/ZxRRqtRJf30wL7C/79lfiXXICXSgCvUBrZBTQ2
WX033pkIuuZMFBWSXJUW/uLvG5QKDPIgN6I0pfdiHbgQVHdksHZCOD4wJt3dTJ2M
OhNsYDnRftiuBbT+mWj1CWoGaJw9CIHmCSYMDnd6lUVzd/eSHK+pDRsgm0yAJiex
TwWv8I43uz6fcApum99xrJtE9LoRl9XAwaW0MIP4wkcwrAjCzPhIsyPxEYNOHVxq
z8DSNkT3pi+lcKkx8hNLto2UgBLYSJN29B2X8ZqFdeGkUuMMszKaZ/SQsfxBGvvl
gnLpZk2bPkhZcINw3zYBRKz0oa0l1XZ+qTMTZHEGAQJwSB7Mm0Q5ixPdDLH9JxOl
K0gjvb2mFDQ71l4NDKhKz84nKOoeZ5FgzLrMZIjOOskWUQ8lC8eNfr9XsVHZqADT
XAy60T1gEUkC8VYHmEA8GTwfPMWMWIqhvkciuPIGr77tWRPfnLZhuOfSONzgJ/gN
cOZlaBP/UjeBXBJDI8YINs0G08urIbZ4Uh6/nxXQiWVWyyYeL1NWLnxKcSTtirES
BgM3m2bG01eQn5DAjJee/a9s92GWLXqlJVGlWGtLm38qriRd73J59uNaP9AXKgb/
9jT9FbxCNC0YbfTVasoJfpo6P/P8iTSOiHMuUuUK5+xRkxHSS8EOpEhYDXS01hpa
3m+nlLhPDR4vVATskNpaYsTbpdFzpLoHEPf24DVg62ztriximUCj8cWEufBp+xKJ
eUqKfyeY/6mkpMBL6+gVusRckHeFkNtRs1NxjgI1wfnxRhkZBeYKRPypgPyqX8k7
TH1SjIE5NGNFB1O5F/PBxi/hlqdhFR5ezmrzF1uom5mqz+jE7xym8G5YIKJ4Bk4v
GgLgZIWEBODAjrD0dl8TfqI88N+DkLWrGKQ2v8QkOFERAsuWuQn3e2/kqF+Gahkr
vdAfsI6gD5+WtK27rLy/M6IaUNkb0Us17wrG29eu7n1XAJlAQfltWscqG0z11HQP
0cba4TIiOvm8sPEEBUWUmS5I+vwZX7xCE1Y6Y+cLWtM3UxO3Va4836XIjfns6GjE
xe9RGRas0q1NYaH3/RoRms2Rhk/XWSC1YYqiprEzIzQZxlobVXIRbaBPzw3FXLmo
gk08i0C3WhlDbDs1ZdLHO/Dcq1i1OtQaOTzmor4rs9lXfK0EazlazgJQ0AXwZ6WV
kJ+2PC5xfbqVHztq+FRJB0kuOiIhomCsb4h7KcUuTioPyMVDhekll2gYTxdEHYcF
JRJmf1vFeLUwXPyp/AouMcqZKhCCfY7QUh+I/urJBgCmCt7qBYGVcIKexG13sr/j
UFVwarxMNFDfKz764dp9dngkSsc7ZaaqasmSQUacyMFNMQaWKxh1DMM22R+8xKIX
kLijrJuaVDQShgCY38fXHCASUZtMN7SLfQMg4UOgtyvMZqKH44SXhyHzjzmzk0lf
lUvB6MO7ie7GaGosxTGEz/A7BD8L33EJ2w9eDdkVMyyWwL5xvax5L+0fmhMA2OKV
hvTFmC8tA1r9XhWf7O9ziXypW5+8w8+yRCgnkzycWmJNDys0xJLmV7By6f1UEDZr
1cXxi6EBwuysoZjPICOiilZzeT5qrZf8zy7dQP/AJBj3S4fru74yKVxn7/dgeITa
HOttrN/PrhGsdInToLB5N2tpgDxpovGX5T3SAZNGx19Xuuc/w5IvqbhJ2/0z1lw/
jTm2IKxgKt31vfbOhJSUxIb/WO4fr8rjLem5trXD+otGJ/lxZgwLLuWLISvjYrUv
g5C8GuxHhmlqa7LpvAq6YVBWavPvKTOtLMs+75yhbUT3z7SHnPfQUb08L3P8YZ5a
27D+3qGn9T3Cg1032++vLoevWKg3rDG4heAOqa92+Cjsmai9xXnwD51qYML63xwY
4b2rUIbdr5YJ+7hBrSHE7n9jmJzYkfLqB1g+XGzrgyGvjRcxrkK2Q4A/cGoJzFOj
VCDgX1pdpQuSt3nmFrSsG7l92J/UaWtD4qTVkVJrevEma3CVdwrgzYoh6OmpdJ3l
FQgPLU26mxiR0TpRsd6seJze9wdBWfKUFFOwpHfthOW3vSDaCzROZR4YGAf0qHzY
d1JSAoJ1NXAlxmE2xLGasgX40pegPehWuqCHNdMtVC4GbZAIdIUhf5e/V0BcLr+g
jwuX2OTgRzOsf2dQzXrd/LLFQdYmwZvebjgK8k+X8+tat3p6lkFfieh3J8pm5jxJ
24maHhzRiwyhkOqzEDSC1mIF8+deSTaa7SxcByj4Tpgu2Wb2IUyfFtNHBcI35vaY
4smzWJ2geVEDkz1NMkngGt3mBCced0+20EH9BQXgaA1U0pqtAqF78UZjQScspwiP
Y9A2cjyq47T0QzOH8MoSB0DZSHWkvEl+ZvN3i3rDujLkriO1YHo5RltCj57TnNXi
YsmUHBddTZawj/ppRyWj3MWxEybZmoYSUF6E+oLftaJpRIJndpEr0ucZ5J6UQzW5
3yDLXWEnvQ2dpgJoxIAW9HRs8s5FCZJHbJbOYX2+3CbB0qG/oyTtSzplHhsT2jyR
J8++E6bHEvSDz8nyyD/srPKnSh7QOEBhxyI8hfWd1FXQrw7gSDsRO7T+9RxV6hzV
VhfLOr9h3yl7WMwiKVLesVR7ItLK8tHllgN4Bhsknmt2/MQp0x9mgMUpUc7HHS1f
xZeul1e4kYwPbRZ3AFSqauHWrt8swIxOlFKllE9gwt58aWI9h+JgeilP3HoVClet
21n/PAmlv+hwvTuBhuu6CvPf6zgD5Yt/RqYzAi4qyICKM8Y8lGYgb2BK8Xv7U9M/
Fii5lumHwnjD/8AyoFaoZUguxWuOi4piTFC7tpLVrbh2qDBqj2HSnCx/gmhJhT7k
MNIobm+gleGjYccmtLNcLxBGMxQZen+VVDGc8B0VU4EfYDh1ptHNtrETb/4OBSw2
LJYke6FNQtektG836qeZy5JvSHyKg3zxj0YdMQyd4uBHTRYFNpWr4zgqLfyHZyuT
QF7w6BDa6wAbnv3VMWn21rlEsMxuLLNUWEh8k4xLm7UGRf9tC4XyL5MES/C3k3gZ
+44f7EFyq4ae3f5W/UW835fXbQbswe5Kw5JCckgAUHpZcZ2ZJW9ds7e3Ato4ePzJ
P29JaHaIhZ3jnKiBHiM8SrK3k6GTJEnF7ug1VDdquF9wkmUHUSF37Bohg/kZjlpQ
tsqRp9uKz5IApyiQofz8KhknxougaL60v/bwnRA6V86xbb0eFnTA6AbNFCLMnFKa
rPtmcYvPkAAytp6IU4bdGBOnkSKmOq23vVJ/HZWuaMbDuxfvEtgQVJhgh3Ghy3vu
qSCLY5qY6uJXzE+fDaIFp5psb55iBmq6q2nDWIa2oDno0mofgEeSOl84XnC6l00Q
bp1flALHz7Dilj56Wl8OOcsbx7Uq26HzSwKeB1F15/ap4jL/PxS+lhuIS4z7xN/j
Co0pBlbbRrQayg58ivYrj3SVMYKaxaVyGkFHjDTSjn7Ua6C03j1J4naEg7Iwwyrl
Kq1oVIEthBZ8fb1WVxmU+4HtesM0Uc/VRQ+/SgAqdVGytqQ4lSZq9JtQL2aPgly/
n2iqbfx3hPPNFeQL5ACEB3kUPcqvyNnSiYxJzS1JkUDZlZO9UyRn1k1fUT0ztFL4
MJTI6kpgUCGo3GJyxd/bLZCyzF+tOociKY4hlL6IG7b7ZiunIeqkkcIoWxJCs+hW
aMa+kYOBC87IE0YhV4Km50rneCJ1y+GHw98DAblR9Lnqaq0Sunjd+JmUudYI0rAI
R5dnanCn5hBoSY1EUmjJWWU2juvqXHfEPr477xWNhaOw8f4yAH582b9h03kyIKOV
HugGUTi6ZG0WsE88aMxMCO9I3Qg8ggqEudZseOgW5kEzTF6xZ6BWBW4DmW0jL4Fd
KTFwyUEhJMp9IHZSFXWGhqdn8SNn9zxnbu9wms0gL7D1zYfiEvYQxzUKuBigRFlN
/nIr+Ouavk/asiH1nXU6N+OPSAD+duLzrQmMb+CISwT/5OZ3eLBS3igYvfxFSgYq
mrs9U6rPvDIxAOwlqZ7Njzo3bJTMoszLAxzHdSjCcqmmIkCEabIJsSEs+XqHphbO
0n+y0WRImMdsG4XNeI2wVX54RFAHFBtV2V5sJlg8JlGE0hrguwq2sDDvBCNvWZB0
bvvmPd4za1sAJtxfuZk0bNTplvxYXJaU2habq187qZHwaixtLI8IkfM49Lln/qi1
mRG8kR0ooNHvLcRcTFXOVvLTJ5ZlVA5mNZRR3SGWS+SynorviFroqwicqm/YQ0Yz
o9Aa78nOTQDTMXuaoxw9jgN4lQXCBEUO83YSrNM6QZDkUItKYLc7kfKStEOCSyGu
jDUpDFAz4Da8fLnR8Ssrh/zHAj56A3UGxKbKUz/UfFoRB2t05UvtX/zBJJYyfMWu
rOV2b+ojUuKs5VPmPQjPYEw3tcv3+A/MO4Yqf1onWVRP7g0H23OJHiu7BQQMNUta
rvUusceP6pAy1FsgY6E+d20tpb8+RpIPrYVosgBHmGmpvl/BrVbaY5sDwU613j8b
zBu/J/6HW3e/rOHXu8EfcN7K0kYeyg14FP2Ud/iDXpk8M7OU7fSnKa0C30tw1s+9
UlKkvO32XrLEAeWKDHmTssrE/lnwaKfarcyAhVwe3OIDcnb7NhilIXyJ3FU/hanq
g0BU4aGXEzot6aJuX2WjNxU3N4geFL35juvLXeke8rFB0ZfzJal56mXFCYZcsbGS
BpNazjd+VmAw2jYHoFP0BxYYjd6NaI4YMr+dej+O/ns9m97gV9rzjqCbixU9VpJI
hy1MGHKBVFpMgG7fEwQZyyxw8yWpsiD67svWjMpzqpCtDVaOVk0U6zgclLzeoPWL
P7kQ2wnoReZ8hWzeAK07B9cmIzf/3CQRKxeGJNKDWt9f76F2D7ZqJSUFvsUG1fuF
BBRn0t07SX4Y8J3co01QlKImfPwl5fELR1rx9j52cK3k37co1xsd1cWbTSy8jXy0
6YqKjts0e2i+i5ri2sXE/0QTU2+uLgEUGfKNXoH65EhYk84KqLZclloPBvyJXfwj
rf0bHu/fQ4OybRrBm5zsL3Bi9GHUDHynAeal+jurGYlYqR71j6OZCU1RhvAahL6u
JjVspRrvTuwRXhGXRrCTVAWAZ/87R1kgMFX/AfY5uRXAlH+Bq3wstgcuFVHyY628
t1Hby3lSSlCezmQgrEFO86u5rB/VdG/SuQ9y+MxKQd435+VCMDchVC3F32vKFTUR
hxjXjIPi0QN3xGOBK/saX3CUbr+Nfl2uJFcQxo4h1vhPYfnKMLKcoXbuTVgtezlW
VWIZkQoA1phTDWorEq7PwxLddP+PnipG+z2tBKSi1+MrKQr0bKguTRKwl7yfzx+h
LDQitqLHrL8LGTxL+6Hlk9mJwjCa7SliCuBeE1cWXNdH3rVuIVF/IyvX4JSFhpAc
LhhsPDMc3YXGaSht+4CvJvKnOFum0FggkyBqFk4fW7X1OWx4Eq3edXUHf9oLQ80p
2Y9w/DzmgBk+NVqRZyNkyxYVt9Dq795L/AzI+jiwTWeyC3EunY44IGHxg7JYrnQA
J04luWimjbUxMgT2WYT5amFldu5d5UxKngaUrqmZawpgojbBc9Sn907+NsmsxdMt
gTNiTt45PtADk6/LpYHzK/kGlU/jIArfYcGKK7QhIS2CNxydVhgtNjNALRHJ95Xu
40fq96F7gBwcH92T3UjwVX5ATa2mguJ0z9omLM+dVw+2CZ+FWBk44JVfQgdU144S
ZWfNfoGiUt5ixcYql5q5PG+zb/QD8pXIZsuHRTpg4xDr9+TKDMwdGYxMlqV/Ukt1
RRuFreSfivbqWD6Ddn9xGdjwmvQ1Z6p6+wjXihGOQp0jXZ9pv4n4aKc2kBVXfNev
I2VCF67GbiWtXw4JySG9nt6t0zpvjP/W8DLAeiRdA63PS5C+e7TMkdA1lnxULije
rxf7uOxgRVsGms8fGWAA0tDX6ecKgSUGlHbiqCWMz9fcInQ6uFpAmAEHLd4SYDYF
rGt04/GST5s4pUVT7+NzkZrNo6M2M387RGSvNgTmq2YsqFMEmar/BDB2X5BdlOa8
wxZTsmsi0UvV18o/nHvuNrph6nEc3eR/VnQoihNlwhsuCEbFxq/F829+pMXx3658
AKkR8+1yKU5TRk17BB9msT3PokzUzewKc/FB9AhQANq3u2hSBr/Rns9S+Eq3D/Rs
8hKBL14GQwnV2dZinkRjpGW/Sh9B3Hv6CohHzKHaSAwmOwAXfcqPCGpS7phRTejG
rNtEQul4HYgcBNIi2uqyAVDVojgda0Xg7MOHiHrBE3IBS3Oi8Qt/dVjN4IT79Pkh
MCpOYBRXMO3fgZUaahETrscGktUpGRKNCt2x55K2zZz/gNSCOE3XHqRF8O75Z2xi
HWfRnVSjw9s9n+vbEE4k18dIiz1KglJXs25QdwcpRtQcF9sD/lZztjgeIWcimWZK
ZQZcHtTs2XYCRJTEiCWiZ4rwovSxEbT9g+ER+p418GUfTcyMjB03cPreETwUd0ML
ulNf9XwGwBSKOwx4MDF4rdHt8zcGZ4L5CoF6c8tTMHO+b7DaeOx+QFiQiYJxte+k
sou2jycyUdMK+pMC11DtuRov++JauK0oUnWD5H2b5MJM9RIvpydCzUiyUiLmu0A5
MP5NipWav4EmtOiNzDEOsP++woWYtIGDbReUlm9HeKtL/Kh4+0wvmo4jIzogF7ri
ZK5F32zneDX82ea47biKgu6R/fOdj43kM8UBcerfu9NO8e7UCf/XRHQSC5q9gWlv
ufZLoIs071q7+TkjZMzLPJtKVNF74ZZfIvj5wxAgKDLZeRvAZ7S4h2YH+nK67P3N
PHxxfgnPAm1jLTHZUOHhnflZIBcf5Dsj//BIBEWtfiJieAoIVg+f7R4FsADV0f/V
SUyUJSYyBfY1mZi+kl0kQ9mHJG3H81zj9PGNf9xa4Z1nqOzs/zwR3Acp7NzF5oBa
Lu0XQUqOh518IWIm2HjGG3xxr77JNSYe/OiEMIPDA7nTptGqfI/AKHQHQwoefD0I
GvMcmfIhtYXFznQfXObsi8osCo8ULNnwZvdvrlDzd7pTzRT+NRHUvZfzTd27R6c3
8OGDlxIhSOCqjsgDCXI9w/Co/HA+F2MdBXa5H9imtvb0zSn8ZW5whVIu1RVNigpX
WEukTYF0bo42n6/z7ltSaX5OohGW0Kcc2WUvIsC8HZokK0e6Ciuz6zldLHm0p18n
khcd8QNjczPvZUG9nUP0x9/CDTwnXB7RiTCczyQXfpeGvZtFuvOU65U75OtRvJu8
KI30e0J4437u7LxvS/EJQDI5UMxgRneZ6+/6bsaU1Il4FNuUkzV64qxB+Oa2bct0
cJcQ+XdUwKxlWKA3txwSWvRmIlgMujqSgmb91vcr65YULlBPq4A6q0We0lYLfmB4
XwUaz7Aviik/GNmE2/96TsVtWvAeur7cSf78ZkRo7CiZgDoKXx1oGgVaFsg87MXh
T0uzsIbwFno/TXhXbhqIOrOfc2jFgF8uO2mFIO3+1Yi76QBptFQIISlk+4Y5qr8j
waNGTfyyCaqEgJcDhXfcg7tJ6l4Umdu7SWy8FmnHYzGzubPWjauLtRPC82xYQUon
/soq7GOEIqnjPJFciCj3yZcPg482LSa0YpI6dpVyOXq6Jv49Dg4n33pLzWZnG3PX
IEHdDWAogOUZUReq6E9PXp+WrnlSLH+xvpTt3RDzIdOqvD38HGdklS3xefziUUOb
kN1CgM0wNVSlw5tULXDQtJBzlJh1fmhHLZCDY8Ny/Vkl0TfczHdvxbw9HCKAFLFT
+dEwFo145bbINfHriXZsICPBdaF9FZUmYkiwvPk5IUqPS2m6zxrVWWJM73/iQXSM
aiQoWsC03gBuQ60ZsVEM58YaU4Ulho0h+C196CduzEavNXOMQSpZbNAwEa3M6/rL
MXPbiPO6CsCPv+qulZKGe7xyel5zGyD/05vComV3AXLW23H2i7WfCo044PS1HD8k
Vlq55ox6S9fqlIUs4YGNSEhXs/CUKsf6IzKs/jMwQZoRWkR/tKOqDzZwG4v6Vd5Y
RXNohyfI3JWlbMch7U3z6gVWcC8MQoJ4/QWCY813Thmt2kuRRfQ1Y3XUr6a16bvG
81smQ+HO38VSGItAKi+jIOYD53VTzIMAhzNXCKvNH4tFwRIqPbOhuEI5aToBoHy6
P8+lknCfeFv3RxQBdRxYzlO+6gIp3jjt/aGzm2/xhRFL9VwsrIrZ5eN04vKddl2Z
ZCMNQIBCe+XMRTTmaTFEGSw/PTGf1fSy0mqPOAsQQGlZVx7Nl2f0mTK4eJiJpMji
WwF0qTVA0J4szccKBJi7uE0oTyPfHQVOw31HU76Y1upAViHhQaEJ9SUD/sm/+Za4
DrHU7Vvx1L2Kuorzx5OY7iju6N+EQ/6S1bYKHrnZbB0+vDinTxhysAi+h1coZreG
dvwHVmAajhwbyoeB8+TudxWnpfCbTNPpvko3vi/D8Nc6BBazcU9maoj8qptiP2gj
vfA0siXvV+usWuyOvxqpdzR8VVIW/S99VJXNkcTaOEYx+GdfkWu3NLCJuqXv+P0T
3pPbQ299I3CpJJboBphN8xZXa4zGzaXdcz+YXuAMsKbK75NNevQW3C0dY5vkpu2a
IqjHFyrsV/rbDJXAGI2OfH92uqlq6BcMPkHnv+qBUUpNKq41m0MFy5MQEd3h3dii
3WmljsclfvPFBuDW4QhLjdF2zZKl7V6k0+VBZJ2msR/0zaUvz2IS+SBgNapTCx/U
XUOc5E74pROMCahl0tmBCYKrY2pYScKMYX94jGsQX4X+Wyr/iCmRM5RAK1bosSbW
CMjD+y2fBCv8so9SfUtsdIX7EpIPh4wx2hpUQXTXwEx7mhtY3Q9TkC6IMA7MboOQ
7/5QGv89PW3xvqVktsj9DKBCYCbr23Bw6afY3ue+zUB3k4ugdwYLRft2huyJsDqc
++NE+jx9lgK7vdGL7XThTdKy7Z80xav/jOOPbZer4xSgZqwwdQU5arfGrWvKawOs
aQlI+OjSHjs4ugtuJhD72HmjeARv2kEdARwA1K7X8jDYEwja/A8xb5O8ExxAlwmz
3ec5drolSIaw1cHezE+iB4z6znJ+o+TXtf2302MTc7a1yqcOZzaVKNbJ4dcUxqxJ
UBQrvu4NhTlNG3Oxa8LRk2EYmmJChyW3iFZ6eWpTGTVsGZBfihn8JDzzWzaQqcOB
LenXMgg6XK5YLyDY9jRFmfq8sAySo8yxIvkBda6zZff94ss4X0jSe7r9EqVy96vx
7xa7RHS8oa2TDH0NiZPH7ORBGqyi2d8ybuc86m1tiUF0EBYIcj4Vh2N2r3lGV1dk
nQ3cuYTuUe4PgQCruI8xXKXnTMK8qM2YQ1mTX3DSfpXVVUeerMN7v+sm0YphA0Ci
H4r7BF4j0MuxgsIZBHXCnz3HPRWjb5ueJrxBq/3VcUWWk1NFX8ZQJb91KeKLjMx5
MBrcXYIvOxYYHvqy3IKMoNrUdz9pYdqws3pURhLk5I5B/EB8G6c2a/36Yx2YwwHT
0wXlpY0iTlZRgHlySsddosn5z4Pks/Y15NKIpWpVc7OywHP6JT2jjBPIVD7AXueG
O2eG2LQ2gOERY3VHXR9C7U+3BB+pPwT+36NjcKj2lWPWNIRFOz7t83LcYoZ/VrXu
SwHCm3iz1MEVjOc0DQTEOTy2x0u9MfiC/+bCiCg7mRJFEfqVjlspoMksvi07zjGw
vOvwK9LsFnXwRQKmAPYT0cYzeIvp0ZofhD+nH3i7wsJ5KedzZgJVCHmLhTBs4+Ju
m90wNnYPcpv21D1Vz4lCAzgWAj9BkA6cy/pyBjuRrj+SSK5tQ4mo99Fjv9lFVXnI
4H+J/4MyThhgsWJiKBdDw0ZUvbuy2q57DeQ+RbqGD4ZbC8oq8b2OZdAaNNKEF5Qs
/WjmJaRtp4Oqw/g98Sf/lKNFIJhmS2IJf9WBRFh20LwzVw2SNFifBQUgODhw0LNx
051y/DcVuAAGRCUHCgvA8I6L3Ci/x0IAs/EQ2C3duGW0tMpTFzhUbkSNc010anPl
trslQ05ZDMgi7JJYkEvB6x1PF3lSipY86QJJvTOBGmji8gdtcSDApqkV9MdDf+AF
MR7IIjxgsyQzuSWRTSBUcSEdc2XeC0Aa6ALn/gdwTnWyOS3Jop62PSeIv9VTRpTa
jNws+Saew5wdOr+6fIKiWscLehMulKp4vr35PGrJOAPhVyXNBWHDK/s0XitIZkSD
dvnMdhtdPkTd55mD9YNbyv17O6MUjISBTTlQ3Rc3KEbTbqh4AfatrNT6Ckm4kikN
rlpZ/vo2pOBwtAeJcGIhwv9da28URie+9ndERZZIxN+6V0dIKo6VLZWXY95rMyJ9
+T2nM/INUF8AhneWe799AgVoa4aa1nfZwLJyK0tUcfgAF8xq51vVKUY1KnhMUsj3
YRLY9P5oMNfAWOkyZYxWDTzm0iKNShUrQGXfDiqITsfg7tSv4rMtQg9E5r3Npwpr
5RZ9YOBj6APvRMth7RbB20y9TD1J2EofvwPwfc21eXmReB1lLUxAaO010pacK/uK
ChrXpAZyS6uQxLUMXGUWLaYyrL/BXIgFH82YGIE1WLdXVT9KamOVIV429jxn3a8L
L1z5nDDX0z+LeMOw6LF1+aOJpy612rtw/pEIkrRGGaAB5bOyOZb7gdfuodtwE3v7
erNL2S2HRSsAdQkqNeOWxFIMbo+Mrl86sA6pXzs6+aa6YkYV5c2JZoO6aURYiloP
cWy1xWqOENrHljFlZeHpOPB93ddaf1+XKahn5R9lJ/0RJaBfxMGwue4LlNp3Ro3H
lTITtn0ilRYyfTP5gBzwAV4EYsgnz14hDSgB2aQFNJfk5nsgTk5HI9V3svrikdmN
G284d4ZSDi+9V2Kj6XyOKZjXcjIQgMydeUVEinhpE78pTQN+ADt0SLqjoxKDnziS
8WqHHzoQ9lKJylLam/k16tZRmB14Duhx9g+lZdMrRELWXF3aDm274g4R3QODmgDL
4XHltRGXxW3lc0cYMdjz+Bmhux+5kiDo0QsRbPnsNdlsqBeI6QHDKGrVRQp5BaNd
dFzQpbl0Qr1uTq/qfjSr0tncIlFgi65hN+urRzQICJJbO4vQOrH3Yw8DZ1UJAVtA
XgCzUK4JZmxEzkhfeEYXLmduW3Jo6Ot79zK4pDgAiWYZI2hyxSs97HLbJyn269wq
+KLtYu25RW2uqVXzN/PcZWcUmFA6YN40GZBdKgsNBxQaGtSGqYoEQnPrd5M2su34
DLAkNkxhJKk4O9Nt92zGYUOT/6x5fm4glimbGQwLC3cjAHkjq/uDqTBIYXpIWQaN
KYzAQPJ05dm4HRtreeh7cM5N6ezoHhBiPjzNZOaJ2wFH9Ux6LRgiwBhawKJ9y2zt
QSni5RokGWs0j6/aXUmX/tragn0obyOQLjyvUyQf8EYJNg8n+98zJgf2irfOiDym
NZBWLpDtFjXCnINd4g3UPuSjDZGFhIqjPud8XKV434uBm2utNfDvGH3ULGPhG+qx
cBJIb75P2ua+6pBebk1FpaoCZhr+gDrzEQpIDt4qwnUf/VewL7l+mZ2id6VjfLFg
bQVJWqXnIK5qmg9vCxLbn9n0bCXYuoSzrcnNTq8Vo6G5hy322ETuG0Kry5DSikb4
ajfPsmOr9hvErxXLGhzTfdFwlILYx1Fq1Yj1lrC+sW/yqOW30zqMuX7p7E4HyJlZ
zJIc3V+B1djIn5tNgQ38juxeo185HrVz+/GvUwti60Jp6ulPE3ar1XJ7gCS368Lj
WUQkItUxcaOJc8erYo9T6OgXw4nX4XJp+oZ5vUNwoGTHvAzpNhofwNQpeHJMVSWf
q6g91pkJGgCtV5Yr0ZUZva8hnuaqP2iSnFKVzD36nlrDcRpOBwUNYZnWNN8HEzGW
72stEbSRMmf8IVOee1YPU3PEkKHWVOwqqwVWQuLXOeOyIDX5nXRYt8wt+Qqog7aN
cVBmxmwwxIQ+NTyYsjTkGoaHnQKx5ZVW+6tvqOAJFtZYXuiMhbfXxWVqdW6p9wjp
UHfdcTx2PYZFTS6KOqSZtjr+midq16rsHN2zX4lXby2puadTIWkmXze9mnRu+vBP
UwTyTbgkh/+mYnwqk3eQhTVE05QNYAGqUgHASNntRSgV34GSw8ws24Av6dTgvgOw
7V0bK5JLm7+XOG9vINJkhWjHE/9VLrBypFrd7YE8t/HQeRo1K85HmfVGg9+edodR
E3Vm4UqnJ78VvJChZYtNHaKr3lL0MiyZuVnbchgVnQPOABmsBZtYXyUwVr7PSklE
vUW2c2wxR8Qu6p/Cp56Df6EURqaPSURvPzACI6vHeWYZ9Snw4Tm6TbQaNmqMyKVH
YMLg7yMrRUzb3jNRFfctG49dxDIOFdY/7zFtev3tEJjL15hWlCmCC8vsvr7V7RUF
1BxrA6m3pLcwX1F31KB2J255+sz2K//RM8+tYpGkVh4UzHNbYzXZIPAOjvxm+NKX
fP3RfpxAmfaf/66Z7cmPak0rYj+3gs9uSeNWkUnu4/g9GAXinEp0mL93zgel2bo2
qYCagF6VVi/CcCYGJFGQBmoKyvs0HksS4L9yxgMGnhPYV+YK9TRzIVwgeCxifWIi
CtyLoodiX8dZDfwVupnP4ior2o0HXwWSSRsMIaO3N5By9r93/siYUdlqeY3u/IXz
3R7RKwlu54ftetKBAPUpUKIfaR2vABT0Y9ccRcq7YQYT7+aWssip/tYz/8P5uE7c
V1xu1nAdThF7gCn6b6PIgxqtDxkXGN9d933KXLpjbklGSKrf3uRjdHq2UHKnvd5V
L4qPe/ztn+ptkSYIMg0B5FdRIly4gt9imeqZX+rWBxxk4DvbfPJnZuDcgUyUAXLI
ClkmZMVbd5YpBON5cjI8J6hqOjWHyLoRnI8vMLxAYg3e6wwLShdLGLz6ywVuCgcq
OUmG/3fDtxxwuFy9Veu6fGMYEqj2eqr2TAxqDHDQBatI2Ojc7F1inYkrTrOxT6Ca
SZHRPzIKOye5eiaY/uCTJd2OybLOMAxB5T5H4ziwSfTgiYMtg7RVx82lVHCKax39
zARscYe3MVDtg5v8XgXLyVeoYLUs7FF5iWPr+EYINRWZstG5WWDodlXbL49aHvbN
XceaVfzi/SIH1Lc4RHMv6y//W5WJDep9p+vVhywMjHqNjZv5SO5P5N0IaFLfLBPH
hRf0gT2swJT7yJCDzaDzMfjNL5bRfgUEYoiBEf+hAXODhLtaHBWvtQTrhamDjDFL
Www/hKFXzhVrQUCZ30zecI4Zl6mMOV4cIjpg57PluqLuuYV+pjShVMsZXXfRye/K
1tj+gJtQnw+81Tc7dsv2BaGFG1gZwwo0JgNYJdr2eBj1QvcbalRasbktQLJ8kOsU
v3qFYqc6G1Nl6d4986wW9VHjGfWw+chIKqE77rFad316dJealhAdbmvy5Z6yLhnN
T0mNdgToWfIDevHoTd07E+w17XujKYN5wHsF5Ct0K04VZUWqxq5Rc/F42fvyTul+
F3dVaLwjFmsp44/RUGTzhwvWcEyGuDYaXIy/JFf3UFwBlgr1y3hLtmfUQcZEK3wp
TagY98B5RhMHADzUu+mcfkLcisaLJdPKsqHUrnSafojP3YGxg8G8CRGpF/vU5lOK
OTDSwpU6S04ddRfcTI86g2fwcN0oZ8nWBx3D+zsoxGvLMklhvDYjye9fjOt2ygBO
u2gmN15LWrb4T46HEJgzFy+/UcGG3DT79/MQJgZ3v/tdxBszp1hTYYt/AIJtn6W0
/01SSKqMLE8ETJTkdf7Y/OagUpka5rYXStLd4LKSETHCTmajRHCchr7+eTM5dkD3
KWreX2CXBrUi96Jlw/W8vI0MxR8MXVaO69jEPWlb4WPQ7vVeFrkJWP/W3e0NR4Kk
dcmXMsCwphFs5ZoYNlIDB4k/6iPzuDQ5HeXfnkLPn38X6YF0FdM5aUIAu70H0g2C
zfTQ79rKKuxJhuZRc6rN4cA2d/HW/OlYu4nmR8ksOdYwxBN4KMZAWdo/UoD5k6Fz
OcO3mNWa1dfRMNJoEr8fpYc93QfYhuU2minYj33GywXahCs3wz70gjQerEaqT8Rv
v1jIIU9oSh/dx/0X+iboP411NisxXjubBgyd3cKfBitsgpBs4F2khWTQGzk7oYeF
r4ZYdh+DN2XrTc8R/YBeqorZeWEi5Nr18aB81HYVKb4QBKnm/m/oVfr8HLDD6C/8
fk9OB97PjIrl0F0U+Vz+3OVWjVikGBhjqvF7k/RBxJ/B2R+dd6Hs5xuQ0n2wgCbU
dpWnisB8etIZIqsL6fJM3k18uJEblCxuCsFR6Cv6aACdYjMyLwkjV9/DSnxDOBYy
VNZ6uRmykyVvHs15dRU4nquoxqoB6D24Evi5Ff1K6ZD7JDX1gRuRnfRzyBiYEG/t
xQkufPzzhVhX5WQWYZdKPfkbB8MchMzNDT8ivIJMNMbXF8YbX1qB8DGSO4j0VJH2
oQPQ4JBJy8j0RMqgaBJarJTD9QrxgHgBQRMl+VBGzF/NtX8o9wDiufHnrhYxYJ5a
HO5BpmhAy69TCs2PdweJJ7i6dRyKIC0FnHGqIswDIwjBjfGgLBNv5ZaUYLR8X/uF
gkU5SYpwG9z83k6EudZAxvkpwVd8xrvsQu7Oy05dd824Lo+L/eprMda29ciQHj7w
+0juAV//Gb9iYdZH8PdW985tFat/infwrvU/wv5KzS/G4swHdc71+wFP+C9AwAwT
JB5DXnaewC/a/NAR08F/OiWo4skTZ+z6nchaE+Da74U6cO247zMMOhGWm4cJxI1i
gK6mMkTJuPJaVHZMWRXsZHJt/x8DXkT4inD6Uznqfql9Y/9Gx5jKo2k5tTSFcizy
+Hx9DlWkrbNEnQYZyr3a8KrKd2YD9Bs2pY93SrxB53CECzGjQhfd1zHwherF3icZ
tvWpkfTjzznaBtroAZpESnvprTm/shadOAfcWj14HQg+2lAHLiAZeOnVKzCDaJPY
yDG/LD2YT7tNNVj99cmYMeOaJVCgTABE+St9+ISfyqfrqlV48kmvMR+A6moxP0oN
L8UBUHxQeHe5qS0+ruN8W7ZbqEoIl3xHCtFJX0umkueRlHN2ZTOyQs2z47Aa25aQ
hzSEuf3bnB7t58MC2MW7snb/1j006qgyxspHc9PgNc6+6jgv0cxX+HUUpX1TQGJ0
YZimhGFLZtWsAyOKvPaO5xkm1ZAZsYkrMDZEniOn3I2pqR3VwemKh33RwlH6mepU
MlhESqybsMlGqhXff4IHJPyPcDEQZACGDJJ1U0wNyBxdJWHUCCnzqKsLguhTTHWE
g0z0MS82dXkxkUroLGKuYwi0FVkUIjx1PR5wHT6gt6iWIGolLv1NkdUzFESaTrHu
256lHmL0YcONemvdP9O0HUki3LWqq2suFg7ibt4zd4mDrA4cc3qgG+RK+373lYLu
Yivw0Kf1YSzz+y+66Q8iMMtAO1weEIcEFS8izi/XbRlOh3rj40auGO2tuMlgtazd
i9LzkLoRGz+nDIgBbgaUoc/NH5LaFmNzM/I+18YnzL3z6TmeJAcy/GhvY4gtUyCW
4tHy3fxkZWwKnYVNZI0OBAKon5mrZYVzHEb3o7FuJY5wpRcc1r/JvSwcBxl0WVEr
t6WDQDX00ymo8P9VaxAK2GXD+sfA9TV7RxK75wSbp0XHbH0m6Y9fyvEjxTEcs62S
lBk183wnYx7RbTJJjoOB1Lq7Up7daV6VBAAZ7aHdu8mZLuHXxR+NMlO+IDDPPJ4k
9HZBdwkH2AqvOsuxOsUjvv51jbVOR5eCJ0d2qs7h9Z3RL4DiJe6RfeWwaH7iL536
8rj75pXWNrL9qXsbM8Q54+E/XvTv7koOL+VPtaDBCG4w00f9aJEuHxOUvZJneFnv
yWnsyRZudnN3eJ8G4C3peCZk1gNL4nrEsRySTqB5CsOACnJCtokWyrYCYMPhMZ4W
XC3xBC0E+On4Wlgav6NiT9Y+WynxEjyD8eobAzE4lZXhd9vgMHv1P+eBH0HRwg/e
p0mBZln4qmT+gYkbWEN6sLCQq2DUFoaVT392VQXC1iksUpECCeKjI1AVNnBe4Cay
h4p9x5hN3BYgHXNIlH3XBTd1n8YwzRWh4rk3imLISo+AnvtbuEoAm9AGhlpFG9Cx
YPkFZDRHT/IGxPFiBdClGNd4IsmUlGnIwfKmEOBuHBiCBSbZt+/LOwb0YxjHeJPG
eN4OBj2Drh/WusoMKnvVFJfzA1q8xl4K2jGKgAK7ffU48+TxJK0gag9Ke46Zo/ZA
WPza3MfhW7SelQ20rMA5BqA3/7F39E1DNsPYpa8CVLJ+LwjwzprzVX8jQsx7ddgC
8Kba5nHdYDUqfq+t3/agYSsQVZacYm9/YOCxdpH/lz+DrkCe4lVRhQGOX2/S/98/
TkC+u3rklG+Bd5hfWvidE7pRkq18PSPGE9q5uyTxNJ8m0emQIf7jU5un+sqqKQQ7
KYViVlCdXo4DaUrK3dbOCdoSj4cRMXv85Mfk4HsTNxMvN5wLI8wBAzkFbstwM/Ac
3hpIE0Ym6dRRNBymhtL7wjXo1EAwlTp4Ga3tAReQrBIIwW0Thxgtl07ldxKN6XzZ
gspmX2vfRBbwAgio3hSJBVw7jBJNsJ0EjsbDhUoTTSjQkmhMp/3Q9GSnQtca4UeK
WV0XxiJxMOBClcM19E0cg8597uI3x2X7UxL69RxwLM7clqLNEPdMMXc5EZ/iwzm9
8VDCUIZ+n/MEEU2K8eERFsqmP+GuaMAiddvDppP4Bafa4Lu+4ciRJP3M65PYsDn4
21PTRxBtY9xkRve23UA9fj1jxga5hvFmuaqvOI5ZdvOfCAvAtFQXXvX4PATYm+L7
kb1j98iGdcI5XodE2nut2Ufj+aYRFVOWuwdiiecl4lGcLpK0RiQCgCja66bixUyA
aO5YzpTugP0Sx5DkMfago0r5U9SVJdA7dedxhcSUTpBUC3Po8aX8ns82YjqIe13z
cl8uwd4ea4DbZFfI7y/r+o84Jd3d2EagQ2ODhuxnlxrIFKvdIGo7S4gBK7V+H0ZE
wsRNo1VmgIhBQN+pQXJCbhspkYIeI12FVxyyVIHM+gJbGU+WLSqVM/ZaXcF8nYR1
XDqBhaKcX2HRGkoBV5uPnM6eY1mLNfHexZYmBdIQsCtRjVLVvv+MHoeu8p0WxJ7H
E1hJY0dgSde7o1hZXTGTYtmyuAbw5h3mPRbnbFbCTz7WUBIZQAnLZjmb3lXVoFi4
0zWs8XM1Sjby9RCbkVkhbOuyPcqABMq+JF6U7qhESobYf1UabKJt2Zxy/RlBSCo7
Cl3rlSltkU7ooPedwIaejwJhXzOU12HwmZhZ6aNEPBR6WmlcFovXOqVfDFmqmhEw
rYENKB+qTi4Yjs3sZKqTsvjQNygxk5pGAsBk9kz9soz7sFcxYynk/amMMAnoiXdg
HHJDR9YHplWsLs16GGyKDJrigOURuyTzvGwLsb6btDWbUXAPG8+nuBO3R/c9Lk9u
FGW0CBr8+38Q/Ytm+BGfASyv7gu2JI9iO5fxQx0ADrlXyfR7O0Yo+zk4OZsCDylA
jTgLMB89/b0y4ehS5m3pnuEUv1hMuZdbKG9Lx9pIt0Fr9VWE9AFyBKYWz9MNqRPk
98gHxxYxk4wiWJYwHu+XwqjMF/KpfPPaB8yFmq+JdwiudTDaVtfb5d9JtbWFb5th
fXY6d7KKHnlYTwvL4ERXd4aSk0TR2ZZQ0XMOkV4BbuUVwI/HtRa+bQjLrUJehPRa
pb/1C8yw31Db9VlYPICr8PPCpRY2tu1j/yhgMk5cHiNlTEq3ZUQV/Rot5R5/6kQ9
vh0eL5xD8u91OYl/tDqFGfyU4oKJ6uID1nmx5h3UdXM7+xRfJDSs7AKmzJLsikkd
dDD1ZxW5vGYrZVaHE8kT3dh75JTQOrxHkKTbgGYao90g5fEYsMzRoQKwUY5FdwRT
u17seqNlxkBkbC+KGQfEcHnw6wUGM26p8n++/J+ru47TQyTdnte7QVJNUuLQNbU5
PshzXFh58+juTZ498zfQCO+r9sjWJ3VZNr2e9j82MHLL+wbFpThWjq3H4xJfKu5L
GOtePiOvq6g4CkkMFQLHVbcPG8vQ3m2KgHeu5CktdEk67z3jSUuIV7Li8g6DY1u8
abAkZPPyuT3s1SKjp2FqOeE5CyhV0+hoWk3a7WFqFj0y7Kj//X3l3jK51AwR0lT5
25qRe/CcXpDvZxL5ugqboKp0nurU9tTeWPHS6fzQucTEWA1Q0DqSIKlF4b3j28yi
DmeB/8Gal6xoF2Bu8sAFfoItAtVxNN+pjwtGkdI1hQHVZ57CzdJqpkks7nB/VHQ1
LInuLNvhHti0lVpE7JlhTPoC+WrklmnBKTSC7t4OypSjvwnwOgeAfAG2O8JICjsF
seDu8G+VLkHOZeSPguLvSJUi4LEGRwBjBM6EVE+WBp+/q/lnetUfzmzmzG05QM+e
OUCfupeKKk6/LCajgUipBSY/9VpDgWU0E2Q7I0impCj/QswmG+KR/vryw46wWox3
Q/mZZEAwh0Ya1rMx8QsfaL6pTgigRIlD8PecqarT2B0X7l2K8tzgUNzGQUMZaOnF
bkgt873bMp0VwqfHfKeoyN3avSjCT2Zvj8YjF+5nXsZ+lNw2BQaYtfVufNG11H8y
+pivn4DgWnFBdkhjx/N6igxrfasuue86gZ098QnwwzIsjeyZUgG3R9fL2AfV8TGd
Dj3qWqLItY7A12JpzoDaU2QdxToYY5HIsAxpOz3v7PG61ezC3XhBCf7zz1icrTMk
lDuln0Cct6ZKj2WTPjpaE9BF+eDONsJ4bS7igcUZgAwTmbjBX5zKWCgdMDxT343R
/G7sIV7b5m6yMc7xlHfOuWxVygwDroIhRE8ieJItQa/OssamZ1/u//veW+NAlxNI
IedhaAWsAHuu4+m6KB9tlmcDQOx5sD1EcE8B3RSyCjVhBXyjQ8euIV2E5xJndYOy
3vKZ7pJaAkN5Y7bvRw2eHvE+UYt6bOUzoJ0OyW5NPW3e7d5E8JGabeKjayGqoB64
wcC0fn8Zs5iywFwDBQ20pdhrAgxK5Xe63glnipxKb92jAqcacJgN0asehC8RFu/U
y42Qq6qADZChpQVShd4Gz01IQvtufPhOWARBvSsowQWTVQa6jLCMwD1sel9FNiQb
jVV+Xzvz8/2pAL6kXenfrF7LTJ6VAU1Iv1rQXevMqGq24aLHJltPEpcVw+HlUN0X
q812BX+zdU7H8kIBSzf+RjFHXUndwjzReYafXYtvwys3wlM9ZWHiynMcUmWViTKI
HEhA1HYXvaTSdZ3udvgs0NDG8cZm2UwyB3Jdrx1MnBUmsOAxIyCKVcKxoYrnrKNO
Gl0p/PV5g5ghfFjTvJ89LJvvXZeGFaoFsnXnq9H8x80GDIasWhe4W5BO7AQ9DcWr
7pGHLx7lSqf0Wh+pk80T9ScqZFCHdyYjAkgCDeM5E1KOKD7jELkJx64bCE4b2dOW
Il44EUYXgzrP9IUZHcDILSSRFvrZcHZroo0liwbKQg48GfL3kIhqyCIm+K4377Rq
njgJYbNP5NWPKMGqlI5KLYZKtoZCq82DQQjzfP19BV2HBxIW1rdcl9CaDVWMwwR4
eGHpI1IJn+yazuUnsGu0lQf35uFFIHXT6esc4Hun50H+TLSoXJLSKtUyar4J9cbq
Hw6AcJfAPMuPgELVtvQAuuGB96geXQNKHm2vMKhD2LONIX4AzcPNubAO/fabJssj
0RRsCjc5Pnzrd2GosaIZQGgfULxVHPHOM2B+lrutR8efRVBArEYxQNRCBppNLiSN
4uWKfgAr3bpw7dJDKRN8jQX1hmbVGbEeyHeve3z9N/v4ruY+Xi/LBARLT2+9TyCI
H4y63IbxZ9QQkSxHbNaEU+2uChBciDYwcs4tw5bjvmwe6AyNHY1NtvT5MJH4O5S0
cR0zUlEzFkROGO6QijDj5sX6sYMTc/1ktSzyWLS85rV+35P/uXzBjrKJfu+TLkDn
cYxujUY4xozFwaJyxZOMYALunvk0gfn+NDi5AjUJ+3lS/bK3HaaSa3sf5w0ONGaa
SSL26yPC2+tndAyqrH1mGr0OYVQJYphPgsOEJqsNH/ghxu5GLsIxaoZOV0uWMBUY
IkfX42yvKJhiFvVmH5mg87V3bgh2EqhQCZC5k5p5EPN+Ak3QT4OGJShM/NSguhYX
JsjH+qUDsRvsxj9Te/ZbpNC4AlW8SFOZm5uXcYzsK3hDqD9n2J+OtdNCVDa+Io6+
2GAcMEGanHCPbHytwveiXYFjX9HC8uFtsJMKls3yopT9xl60IXn5TtUEwDQctVqu
y/lZO3K+e9uFhpaxstFmpr2gj9Oa84bkf2tDgV9FGINrciQYGumITZjPGqJdiMkn
dkyhbRh0x68ER1uE+f4nncBzFR6O89bHTJf4T5FVgQjje2Ip7ta1EbW1SoLOEeSq
ofXZ3sDp7GhgVLbbiPAbhi9lCRExwphvJ71sU31fBmaJaY9IyOfcPiJ1ERnrjKqF
GGXlNWmXG0P4kBeIfcu7w7XjoP/7klqXbO1M9M/2rDbOTmFkKyrH/r0PFGYon+pc
mLKeRMB3Ym4bR/8Pw6EKRHGv2BaSzIjPhLMqOFRmKGKJjAtfSWirKSLnk+UGc3Xi
RQfhUDpaMaffmyKAz96Lw5/y0ulLR11QuFpoxOTr1e/KuyAUpI2Xkd/SMbfG7SQD
mc68ryf8E9bHkfuiuyuKDP/cgmeiP42ejaWWOMIE0QbWRSWcQ3vikLd2rWoFgySf
jz0Lq7r/f+QDSBq0FFfPqtgEnLhNT8oEy2GAuONBEW9Hg+07kZFByygEfAc2qwtX
A3pC7LvCKUY4vN4x4vyiBSjBaPdExOCIycviv4XGKKvxhNKWcH5eeFWyrfYpg4w6
kgIO8rDSdrn4R30tSrsFUWMy+PRlbW1pYudHg8pI19a4Tq/JcG9ZPxxBwLKaqeBL
ISaWrKJgkGjAYIuO07eACUhFiV+6oVql+T3+0SlyVXF2K5SeczlnEBMh4PL5yLxN
yEPgF0f8d0MaNcgWEI+uFO5pg64hPKohdKTqb/5HdvD6VUYkizgGXfl06pN2ZOWo
8AuBTcj62A5q2eR4bZnO2/u4kuAWlVpFsEnKkUpGcTnDrXfkVIxmzSTve1A28VGm
q4nhBt/x5EaOYh8MTpqhjsjncnWiJB7jP2Taq2Xfk4qpGVK5D+C2hhgECYUkYy3n
C7Hkv9Z01r1zOKNF4NcVKRBi4aIgnnHKPGnpgneBwd/Lg0U6wWxWWlsB/yJEllXT
WGbdaEvPr8ZdCgrpwgRP9moqdz7T1AjuqNTIdFXABX3E8TJduEpCrY0dw4/xZOI3
h9SGtyYHEbeUuYuOkfwB+xCuw2NCDiF/G79KZEx7eA9OdalCorm7N3xE19d8Bm4A
ayveYIr71f7S57D5Y9rufgKf09M5S32S0Imi+ZZI/Y6tLWJ8VG89R+nmSpLFBN2u
11Sfr2UdvgAnYyozyGpMHdZ82LS/1dIVvdyi7rb0thi+RSHq3olOGPN/MG0WAvoE
6FM6CewnOI8ZoqxrVY4QspE3+5Tv71fs82ZZvUWrX18IhFHXeyGTQ0hEMwdnxuHl
2SHd5UxsCtDwGoAd9EnqQGIDkcEGhs2kGTR8TUJ2hA/98vejo0HmWeMBf3Nmw+4z
3D/0UfTsqyBKnrU9KIeHKfRcPeZDeLKHefDTQ5+Yc4bYnp6SJKGn9nXBp67+0gye
j5SFhv/sMYSlWZ8voDmOxH//NB3JCCa1/ljJopbMBd5eBVBBUQ6mHBb3X+nPWQxy
89iQENCRWiRjQadu5P5fw1ruwTnSkb5vifRiSfe3N3iAxpAtD3uhQLBb4q728E18
CnZ5B6CHNZNUnHUN0GeEZIhguOm/Z3EUCdkZq/11T8ecrG/hvUI0RNtzWgahasRC
6rcW8YbXMAt5K9TpbRSe7+BzZSt+Khb1mh/gZF8nKhPnPvrsN+rpM3zYQ2qGTh0r
sBOXeEHlOzLVzTIhqypTnGX2MydufBcLw8WE45hHGdxdruSOFF/Yoqbrl1DZXuCh
NRSKphS+MCB/ORNtoEislRsCYn98B8hr9B2Di4yGjxIK+lK6TKvjRxfa0j3fu3FF
GV1VLdnTO73OOWoYoUkKniAuAwkAMlcTBIc4urwJ5sfAYRpGDrGz14v0yjdT/joU
FzphO7BDP4cpVyMFiyJ9Ru63+WTtZrH5PXyz/mgTWzbrHkOY13YCOY+SdEtdrVoZ
6X+18juvAk4yOuNUvcyG3eKWBdFSYArpT/EJOBLbsvBOmXS/pof85Z0VpjwbMl/d
ZC7bb6wL3gZS7S5b8x9AxnPOnkgM1IyZtqKG+7b0hCn8dpAQ8R4Xk2JQFlpOG3Q1
hRWgoVyrdEL5CxUT4/MPCxkOs43AOd92Jm35UK+VqZ4vYNyJTxBSQ8RxGR/iXwBX
6Y/aZxwO8Z/k1HlRtqVNko4gGHQ/ga+rz321YG3Tn+1512CuQtd1XhV/GPvD4oBn
4+Wf9gdY/eLOORkhjhVbBB1wMnCNYYbtnBXjooavSxxBYHEnwpBNFTvedEqvN8uJ
u6lbfKDEgdjuGjnP189W7UTArNQDS192rKuBSyUMYRee54k0QkAl8fx0h80yYQzl
4MCjZ9ZnKtZf58c30knvxfsy+4THAslc4X6Rbzxb4QVCWdm9V7u2AQLAFsNsQV6n
ITQR4iSYU+VEedsOjdTSVHnl9FiwHKaODspt06UaHtb0stQIOSv1L/MtBHIXQjAW
I27191eaMpLQZroT4iMbfPSbwaxyeRVsCu1D/Ow3xAhQAIgVURs72qi5LfCpYzec
v+pJVEpuhfj2z1Hc7eU3OKGXrHTpkF4l1rQXCGcOCcj5PCiNa3IGvPbd0yWGuHQ/
Deaf4OmLQ8Q0O3tUdxvxZ0eScHxgcNkbsmhdrlND8bvlbODJvi5seSizWVH2V3Q5
zB4PzfWcdzWsBhY//uPpyCBznRUc+CsfMCXyPJpEunH28d+cGP3XmK8hqsg3TMl0
lXTEdu5PSmomRCfcL6WyJ+n/QGvYyA4PV5Bqr0YNC6fx9CaeZPAJEo3hTFNQaAaY
pe7D15DRE/mfoI+H/4nz4dYBhBrGu+Sy1GrOvCE4fuRsUVoVxayDTSSbX0P03KXB
z2ifrHWOojT/NSxXl4KIdVEsgvprYwjh0R19PD6mkrq9zw8zQMqs0ascZrUWeHaU
5ebd3Ug+biVc4X7tGEJZHn/U3lS25iXAWM55gZmto0alT5d2uwVYEmxcTsrpenNw
5GTEzc6bBXNmGEIM8sxmd+LegLCZNs1F++SpmGgHFiMIhwdRHUo3qjwMFbZetEB2
uZJtW+edUASPmGl4aEi5vRIhy/HtUuip6FIL5DOoCAa7dWWK6nSRkGACNHZwXWDW
qm8bi8r8irAjpf6pVIgg9fYy3ieh3B0iY9WzRBdKgrEcrYKIXPf53JnLVN1bbUfB
IbdYVsp30XZgg2mmYS+Fujd4jVnuZF16qFA8rxlcl+2ZJG03Qm/jMUsPLLofN/jS
b4JI5qz+Z6LzIhFxrbgHQK30HcoqgAYGXVlA0+UL49YDITdQAQLKAFkg7oOybFh5
/PVmK1/5x/LY2Bnpmy6lNJWFQC48naGe3xOQYIrrMtuyoLsXqBmCDsZPY2Lb2JkM
+14Kw1iQwuDNWsmqKaWYK5sZSDuvUbbUbOZAX3LBpNbYe08yp+Vm3LbKSUpAOUUM
qh6T68x1fToxaTSu/7GHxeQLiCcr2hE2y5pIJrcJv0x01UQ0wRF/AaOp6qUv96LR
mc7PJkqatzi8LHWcNt8/hwWHceSoLeJiDLGyB+iaF4Za9kKJ+Yv72sf+9HJeHPDn
huRAwZIWzDN3L7W4ZvKrg02nycai80CemcOWJe9RqAt6+9+1je1RZ6pNGJDiC3Or
HOjmU8Wr09ktLft/xebyO5WfE0L1jxcLIejZ7vxRybzAx10LKwuhajoaCQMHt++1
ma/kxR9mAZJXlV+hrsxqdUW639SXLd2mUoPU2e2saFgU2Qony8Afzm7zKk8PvfvN
qiKZE7AwNJGbF5pJEjgFPzJnU+zUAahwbdy+79xsx5wrxwiinopHfHlEUY7wenqa
Gl0vrWTzb+bqeuiZw7H0qyza95O79b5KqO89ZaFq7fq/7QpuNPvSAmFP2tj+y9NJ
75Qkn2WGXNLndtGuaLAmOgW3M3+ZLDH4H2WdTqyLzI/yZqCoZIOXUyJ2UNsWrBZT
Egk+3zJRtKZvI/uCkT7y+BzKWVd0lRqSl/AmgW3NxNjDW0SFTGlgY4mWJRRGRtne
A3fCNRaRNjl5tMAK+wpPrzw8F0RHVx4Hsuwg7uT5li/jSmpnX5AozPaOZrXY6nJw
TaVrCg4KKeTRWjkQPyaGs+NZCcrh9bEvmZvWsyXlO5t38gzaJ30hCj3nqyfLgq34
Hvp5ixPBg5wAEaMMsGcF7jPDastQO10kUnpMLdwtHatO8s3iLOjxBH9G9kpJV7pQ
HjqUZLktoqaUEmBk2K9LrRSZrZEzySQL9CcW1CCG/GKbROlNXBLhOjj4555efsBa
QNYj+JNZoY1K2V/XJxiPmQxjjkelpCGeJr/Fvon9fb6jvRUUfOFzK5OtGoZd65mZ
zByXHFPx5/1YWK/xMrgrMnXTw0to2Qdm63dPe2Yb3mZfd9Gh9aMUw7J8b9xYsHjq
sE2ICVvG3b3TgEGGZiGqkoOLjst5NNgNDtuYUOo/ApQmb4QGiHuZUd+CBMzJx5HO
K7dsPKTJZzlyaBKb3P7mRJZC0NqjOiS20zKlgjomA3vcPU1U8Ly9ZCPy5O0Vt+ul
orTVY9zzi3+HacHoTKQKBodTmGvXd9NvSrCSoMTMfiLzkK6xtS0PuA1Q+1nSAB+5
Y5C6MgpJI3pIgZoNKCr6AQi845Wucq55bI4kYsDao5BQH+5yW+22ukhsl7q9j6/q
nSCuS716w3O0kFtaOCIW23zuGJoH7gd7oJCilCMmPwLRin3qHOtQzAKDbSMkMAvw
I/pHLC6GHX2z78AXT5IYmL4cAvVDlzZONvJIsHROIJmQwyCcQ3uyipBnShIzDzD2
0kVHxsbh6eEvff/dx8G0D4pM1JPZKBzVL8agGnbBnbcrjB4EijbXGABAJpOeqUMN
PbgJANxqnPEb1Fb04HteTN7GeXghbB2lVMbXlnXEOZIeDwZiH7usAK7AaaiM5Q1w
c/FAk14CZ6dZYQCPBw06jfPLi9cMjFzYWfhpi7FjpnkAclA4DHJN32VLbQ3pHVC/
IOejw7rAb1CjfWq4S2HzimUqp5ybzGqmSaoIrc0Uzs5WdZiKRMCtpCYXPYfkE5ty
ARM69lz9LlyDCdLHD1PeaKA75Aao8G1ZxWLLNEDcvv6mv5Q+dwZWJxTZi6yy6/hH
N+72umg32dCPanjO5JWCndKpI1tf1nuYtOuolEtj15Xur45UxXztk6D4fzGvMebq
n3aWj03LNTYf+RjZ0ola9simKCe3D3jAyDgW4wcFtjbCQMxxY3+eV5KZWiy2KMJO
wWRPXJwP+zgS+PHLJa9aAjcaAlsHSDSPDicAAkL3Ga9pfeWG2xoX9N+gOQr24Klz
ikVwtGvMQEXz4Qbv9A1022JTYE4IHLkPcReI3wWzMd7RtPunB9Q5TEZUnZhUST7U
4TWCiXh7GnypBwpZwRnurEb/XbqvbTGpe09arzKShC8Avjjbew8SL8uIkMp2InKO
15bY1i+X4eRmGqggNxTrerrD7xOMScpfOCH/K4Y1eAopxJdYLZ3k2Ftragr6/ZFm
ueDdARYfbBvwSnodySV4DrPhsVdANPenwWYgAJld7mzWpEAbF9kiyyoPuC5obeRz
Yc11WkcD2prCtXHRwKbvR36hI28uJ1mxLrO0gLGfm2lk/nuNj4jHEYM+ZBXdHmbE
ehksjDQ50tEXOsPB1U64Wod0CfYyzN6nZom2kDd+Dg5Yuewtm6VQ/QQ3SLWx0Pyg
r9jSaGWMZdgvvdzoOXeyhXNux4Au29/46A/qxIGuf5HqAK3W0Ew4PQFopEP6I9x9
Bc+Mwvuisn+znHVnEZCfi0xyzmevRvVqD5kePjIEvezkBl4AcCeVuGKBwF8617uM
uf096Fb5+XovuspHcThSDqPXo5lCWXKTt0Xs12v/OqjPGDi4cLYJuqKf5z3VGQB6
y5w5jl37MEF/7DqY9X9szcFNKwX8rOVl1rW6qteeQ7iIOfeLMMg9cVdk59SQ2FaC
Qo3qCdOcsgEicNxPlujJSBSMEMjSW5MXYfLV+f/L+cpjDN/Y9aQfnDsV1MQywUjj
uetiFJX6lOvDF6wwaD0/Xpbip559dYB9hHj+EwiC/dfb7r2TwME0B+DGvUqpGwwK
7V+FKHIi0xLX2uZRlF6MxwXMDfLCZeJdKPTIOFGU1O0eWtMRK579yq4skoOHe+u2
/XOLjeShdhDTAHBLu4DBQ3utU1samURDWp9cQtDcqvEC0NYCv0SVm068pv7ubMZE
iKOzxiotLLuiFolwYpIG5XO3dcZvflpvoguMJxrfHGvJl1EKcWv9rjtrp2BxEMr+
V5U+hd9M5OIMmwfMo01r7toWo5kmISJh2RDap9mFhZxQsEUnzzwOsWjvdpZoqr8R
rmrfazTWEGhb2uw0e07KNop5nnq8z29Nb43f9UcBHQRz76vFtDUlASRiPt9khy+9
B7fNrXxW4uilS/x4bBfEEZJh9gLXL7tP0NCUnT+qXc416eHKQNOE9FBHkDG3FBjd
bK0fbIZJrss38fRiChDhKGjO6g/26p9LJpNsmxHe1EucauHkp8yK/g5ALcZ1K7k0
l+13cnKgp7Q7t+vgCNV4EGlVQ+aaPp3uaKOgCFmM4M9SHW566F0ZcM3m/jizvKkH
BFNyELYRPs4jc4jFEYF+qHDLmnnypAzG++PHO3KlolxMeAjYjAnZmR/i1KeaXCcw
HiTO2GCrjNV1Rp2sBln8wVzlt4/ghMZPzpXZF+O/wJreVA+Tv+PpPmLyNhLBnVz1
mDMSJHVbsbrXN31dhWmiKTf0JX2RZeyYYtm2eF1mmVlWwj1tO6cnVr3U4tDXjGLG
6eoJH5sq8aEC6RCdNgIGTq/S+qiXi5FACYiEpCTFsB86ZVGNTkbhGitnNUd0kD05
QFLoQq4hAZdBePVRZi/Y4KEriLhzbZ9XGlHpYYDl9a/fx8mWphT0RSxC6WRS8GVA
DBXgTMC8QZ28V+nfw7UUCxik7l4GGk4z/UgWw+qxoPN5tZu6rjIcXa3JdcM0v9lX
UE52z2U7wvt9Jf5dC+cjfU0fW+cFQDUoIQocJrLmMkq/R1acRZw1ykGr3HCkli+6
8/HEVANh+dmHa05EsZ3oR+wbJsnsRfFoOoP4qqSvdE3v25+a9eYXh2bk6iWJkEXS
spOHrnvRFOUWZDjL5qgGBGAH9Li/5IZfdCm3CjpF71UUB+lcmiZl6R1ByTXqO2IE
ujw8EBrC+xhkUvk0Uj/l20h61a/d0/cdsoJuyMZOEfPMJEFTyZD1zU60Td9OaIJx
upKv4t54h/lw/Ho5bhlTRwH1S/DG4KOoLGRdBGW9p9FPDIrkXxPjsjVHC3x0+xq+
vPq8ywrwwqQCoJ6dxMCmZ2Qg3W/3UaSj/TBAozBQfrEkGxcIdYiz3uDLGIEEVVrS
wWLXoTbiydHdg3bTowrG8cMudsgdNNOxF4TcmWFrkmHwQv/cdDxmsY/wGfAymLPx
i/yKfVEiaton8Jt6B0P9HQMJMAF6aBscPdFfcZklf/kEYS+v7jDaEYKK4N6eW14f
ZErtqwj6lWukX3nF+I+VUCQA+6kNn6DUX+rvIfKU1/N+g1K/Bp8MALCMbSB07IcX
3jsKnP39lmVMRxuXkrMHKhwYWQgI36A7RBxB6yyKKcvam+xVgQ9ls18McfsJ8wX2
4in2wPezBLtIMvoo0WstUZq2JIQicDjFKwTqTsjTKn6JUydvJ6VyocGMV+VtPEnk
KkS27msZzqDhJX0N7KmYa0IwKK6pYJJk6H9A4ldhFyJ8FB8nP0zYqQnwtqAMci0B
e2IKSY3HlSLaFpTl2Ojyh91dcSZKYQhanJOW6CKr7BmSKOe9oTMdwundOgICgpqi
75PYlwocF0vaGzxVSM+D9BXYprCZK8b/0EWf3wi8LI4oFVpebCLPte8B9ECN9c7R
BT2uVHBbX/j8NspCHA+QY29D+56JF05f9GQVt99PkK/E5nXT26N1aJW4jjsD8JAW
5a5iYyig5z6qA3XjHP5gza6fibN42A4Fz6drN0BNM44LMspop+HLF3e9orpWgQrp
NXF4FYtyRTkk5B+TNB6o2gFOl4Fb3CUM9fpn9oLTP1mervVUPABaWMSnhgn5lUKK
irfy/8O2oeP2B020BBt2bLUSlzvYhNdrBT3Fx/Q4SF7bZ+f9ezw/PzBIp2jWcn78
gAOpQ9DwXfb+cnfkDCJ60dfWc9JeYbSX4iXKOxI6LwteG2Isjqs/5Pk3t+bilGCv
Luy8pbSkbYVhz7XNRQuEHOMh5NpDSsv4DH0e1Gg0Y2CptfvfFZw6XobovuiKGPdN
ADgeAry9DSJxPhd2RmZ3TlkwIgo+sERe0fKdDIkJA75eR9sFXTw+zsbFY0uymmss
Qu8tDvXKsG/ePHKiSwjeRoGwlPZNCO4G+tkAKoZRQ5G/vbg+lVQo45/3tPP/ykuF
D0op62WFa5ofBJy2PSg5W7os+BYBbaGKvXMqBpXUxHxoTYlkFj8cj6L3tjOyAxEc
43VpRqNlwLq9Is1NO2VlqZPOplu6B54ElM5Oxax1JeU=
`pragma protect end_protected
