// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:35 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MkHvH6FynKlKUqoF06/8Nb82ax/MvRruT/1PqFI08t5uJoedOsbYFZ7p8wzq+tRU
6kJ9kiVjsUwurmo4f/jOE4Pk6NUzfzAC6/UxBgjLfxIfU6sua6/gkk6EOyqXI+Mt
M36g8blkaYAzlH0JhG4S/Ndlb7j5dA556c5wsrx9CO4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5744)
DUM+oxzt1u9CB1EamDPwiDbzmGqzGQXLhrTbaOznyoVeEWhUq3uM5vGd8ljtbYr7
e0NaqDZHSHhVIFQMO5icSZGcbSDF+QezGNm+GaawNaKnYpzEHOLrHsTtfTxoOAGK
5/xI6Sk14vCu/7D+YVhiJOAiWqnkPTnkqbvLfyXA2ceCwCDZ+yiLUuQErC7dbKVk
ght8Z+M3gs1zKJTDnmjsx375gCqR1aUVUC7cbxwR9G9Qchd8htXoeeCWHxMC3Ojt
5gjPKJhfW/mu4s/1Ufn4TcZuigu5DN6A1avebFeJ4oM5TPL2BIx/yX3wxFFFwMB3
cdJvT7yVUHos0cUV8+y2mzWn/Kgtxta1JZjVSgHJVmHP8lE5wpNqzKOzhgJ/jtEq
BTto6OX+v+pDu2YJAZdSwjEjTn4rSEd96RZB4BJvY4u0lAYN62YrciIAwKwIQ19f
vavl2zlhxkJH89FO6EPgOA0C0pqeTwWbQ5+Z+bCT++iOaEtXtiRs1iEPhD/DBsHx
rgH7ZZ1oqKAMghkFfGdbWWwvgKqb9y/5uNuqC5+Lo0w06oT/8ACCRj/2jWKO98fT
TXsB1Z5vtH7exOGVeZJN6P6azwv9234wVg3uGbFRgSWkXNr4Z+Hz9uUPGqasXsA8
TFygFBl+UGenB7iGHJh40fz1GODCHkA9lIkiTHX5QkQ2imq/AcewK0iRFShAt4Ni
J8AL6cnBd/yHJaSSXp2zGnM+FTpO4258QiQ6j2tby/uP2ac59p+l1opzszzzIz5p
818k+4zkn37AeB2Mf+O3XcwDdR7339TtOng8egqN9EihlD2EUX4AKHhxYjEixlvG
zyt3lxxqPMmHNX42KXEfp10oegpgvBkVpSfUZUyjHkMS5NUOrKROZc7s03+3QkaV
WXCx6jkcZ+X1tIO3DfzPEt/yVlfdZsjoAfHMADLT6mRjgQGgHfiXDbxxFN2jA8G9
NieLon9fc9dnmCpVeuX3UWnA/HES4qE1SCOHahaxFoR+JBiSl3YBKwq2XcFUm28X
NR6jcmtXtnr8x5hu6SR8E7tf98I78FfJWspwEsaqagXKj4PXmykJfxHUtTDm6Tn2
RK9EXltwBzQtfQpg8z1nfissbD+l7pYYVQf6gc8Zf/g7pdNC1/dCRmxnl8eXkuIP
6Wk/Zn90Om9k2Utj4HyNRaxRYxP+Ddr8MYjaHHKthoIgAfckdJ2UZCVkziKLBv4g
+qHRlGs0FcB3jZfM2yFHhkPtI/nN7klIvxbzPXT0u1lex6eCIdh4dB5YXfwdq7E2
hfjJf0YQrCoMo5esWGtP50rBuhPL3j00INmV8Bz4jImqNyu0Q0XwhuPMF0qHLSFE
dEu4LxzX7Nb93CgRiorfl72s27rh6uNFSKEvHiiZ9G3a7MYEyBV3tYKer38sCuGR
1zIgI0vpl6S7DrKzwr4qK+QB8nop9MCTWBuLz0SNk5Rb9KGZrykX5z7URtH4OFEr
3w/rKXQsS7S3myGRxz2wZuwsWPpeFqAcFshRko9JGBtXUEoe9IA9ZMRcEyU0owVc
year3aZMyrk/2y0RFnZNDmsCOuwPtxecIbk/GVdWnQnNz/GThEoGlKm6DfYC2QM9
jl3BCo2s3ZgWAOSmCJqf6KrFkqk8Hq/Je1V7rYejuO23EMNV2PB07w0wj4LIpvse
+fE+G536KSlcddnbRWsiCsJ4PyZcCQ8h6J1GEKNzjB8yDLDJ6b5aRp0PHLML+REL
T6ueakJPm2S5gfeEiRnwpp4sm4SdaF+Wr1Q/hbFp9iZR8//pi1hF2Q4n4YHp/dEE
KVOADqNInkGzzkjakLtRxJVBlbe1L8inHdH55GZNWHUKkmpL2eVoaMC+mXqef2Ib
lrBo47iHY9eSECGXEAxz0XDLHfeLlU1aP+c/8CMtFXuXGwee4DMvZl71h3SMDAG1
+R/ZW910kPce1UUeF5IC5iGnfz9wNMUXqlc1GZ5Otu90d1o74bBUWJlgnSPg/0NI
2sW2+19dhpNG/4UreEStUJ4hUWvlOGWR+aNkeYtU8tLLCsnP9MylveNYZeXdkXgq
gZnqgt5e6YOottMnY3Rg8BdqQKChETviteAtcHIdvAE5EmiJ4I8gnJLty0tDAVYV
b5pHAq/ZaO2ACCXAGFmGiv910jKVFgRjsCkxQjQZvLG4rrafYu1y4iQ6d33GGMw1
hzLWk1fUqH4mMuYfMFtIhp4V1iBUUnweUo6/JAOm8gFp6gh95AcaG21JD1S5ohSy
K/4XOdD2hwItzH4J5UTDCnJ8vGJQBOnAwmj/yK/YK48Qq/Z9uN/YxBF95cK+IDwZ
JSVtOjsGkVu8oMFLnxMGiIq8yxLVppDOWxkb9R5QzBovKdTCzoFc6svKh4A9/iQi
O9Yr1Et9oITbRtCTqI76hqi5GANt+rOT2a+lHJLBK7LjpR3kypmErptyJys2CYEr
31yscaC3e06pmla14fJ6mLY3Fj/yRT9FVk01QFUS/rtleLL6BX2yVzXU38njLDZ4
QVKurT8sR7zBOiV07Cn+pzZH1PmboMZ3t20uSXab/Shx+gjULYiVwKLHwdc5iiNA
+7ZIJCbPRMLjeGQRZcIeDtOGU3f8nkhr0v3BqKRT1+N7vyw1qLEJK/OVSri17ZwK
G2wxIdgR/8rSsgjioCgVPLpYJeOdmqsnwKQrTvTTZyJeSQEVpNBhzpr9Rr1dup58
szE+pQ5rQ1xsCYdwbYNZN/UbKjwlmuu0mjM3GhgX0dZ6uwUUk6qKhw/8HgHk+Uqg
3R08fQ7lVr13oU8aSEj2PO2j5KqyG/fcdzIr8gJ15cybH56ai54TRVbhdi8yvmz2
rxGF2ewMGYKItaevmAp2yu+J+MQp3oDYWE/rpN4TuRJ2C1q+gHChx4noQe4g/FO6
LiguWw8seROepzWtPnKammd8R4yzXWbZftlru3I8C//7tM+9zwO9BbKNohIbWTCi
yEDXv3ND+xlBdXVbp6/CW9gxyuuvlHR0+f57Yt30DjyqxgeNhW7w1nomllunKZuL
rPgrIVGXVddo3x4Bi84a+9fEHXoecjqgejNezDlLtspNtztVQgqv35oIS1e2riOR
tEd+hdJFl07U1TPfoOHLATk8KeFPxlztp5NbskvKE9Oiz0crZxfx1lZ3iJ8Fxe15
pvew3uDzshZaC4slMbxSBiDFTqsX0TEu6BUec03pvN83Qf8EsuKM0pZTjKmRl2Px
eKry3Ulf0absKqzh5hnVzSqlHrhLFvmVAXdjW6oYTBSZBXrbzXDFn9GI9/8VPQOA
ccDYye9T2T9D0Ywony0S/+v07AXY186Lm/MKCoNL0cLBI5O0VPaqeKOERQk5bF+h
m9BCnSbhfbIwGH/LfG5V+vkd1MR9GVCMpCZNVxwMrAbzqWN4CP7bcfr3EF/Hy6+I
V6YQClgsufOIztU1pa/LhLEpcpAvaLQucNJXDNEDeL/moWFSZSo5aYT7gMxeb7BY
ocDidMeJLcRssXhBa3oQqM6hVWcMfmOSYFBdXEfuIhHP+pJoUxV1+i5Z+jG4fv4x
wfc0p3iLJufEeY3SfwDVdtl38/D+/+p5AVcfNFWqv2Ee/HRX/r+JWtprSke6fo3L
L3677V7z1ic9GUWbQ/PxrhSDFmwSAG48P+OMWX+tnpS38I/111O4LxkC3FF7Qo2N
EIFLgCkVkfwzMSrAp6RVq+eFqmebl23UVz2+XTTCW4dAudcFSSNh4Tft/FFsjLAf
tM6zSZFmB9BnoXCBRV1+/esqUqiA/Rv5EsMd667bE6hWe8Ctr48iGXiois5Dom8y
+g+YkUa9IKZkDjHI2IzwVe4DtcrfieQVSLq+8BptEso83yiF46iO1RBeQlw4eUPu
UO/HsJ0FfmPhB2sYuZS2m3c0jwO7JErJodOBh4sGJsCO0LFxj9vpnV15oKsCeUPd
3nVRkFs+7gAfnAbwm9k87iiO9ZNTqPle0HWa6h+KjnZLafVr4q6Khi8QNXBEhzyq
hrzTHRyLWDnH/tl5fLHZeRCUE5nmPnWw9Y9MGndUylgRAN0fnmYT7O/pHxhL8/zp
AWU2AwrDn+qbIGydtOIWiQ/AOTaYjDc9uGuzkjfvQMDIgb/pvWnk4xUqc39xMrv1
6dcKXkI6u8QwFQ0+QHraP+AF+WUVJ/RsKBzvhDu0KKcDA9se7vnKEJ/ziwQ9Lvd9
RMTRgtLuCAUDyrBlu6EmUbXD6QW9ZedmEwrCT4R5s7lRMCK6aH7s1TFqCMw0pgIG
A1WbcYWMZEgeC+Uab5c88NDakgmpg+/jSuscz8E+vWp0sqDQxysh9ZCN2w+FFZ72
qaScjvWm3a+yqcMRQYxLyi79B+tGu+4+BSG33weiRoiw43CWsfHflVCDZgy+Y1XD
YyCKSQPjlnHUxuH3rGVJdAkWhCWizDaK8qzi1hvEMjsuJL0toiX/ko7tWjBsdA54
lq+XhRmGIk6mFdANgxkf2pjpNv8z/ezSHjszFpQP8HlovoRzXM5pS6Rkd+jGDmaY
CTNCDLA04N/qP9HMs5kIVhaTPj5abytgUhb2gnnGoeCHEKomueMAVqgLYPBMIaFy
Sq+qr9LYIE9NvLcavN5RKq0bQ6KjKpSp1OmbBsIuVps0Zgt9CVS90bcBxjGrPI7z
ThYgqLcRxW7NgAp0/REPrKmSbK4MCrvDW3DlDc4hHqd2X2rYBtaE4Td65p2/G8Va
MAqgLoSckvzorfWWb9hv8vD02Q7sSCYttTPnYlZQjYh9Z1mOiustrHPMJy1di6Pt
iGhA1yA9btB+4LVQ8JaPWZZJQaaJ/M2hG4oWV4+QR4L5REt900ck0vuCxIO+y8oY
O67gmURTfMKvxpoBvUf41e54qzC+97XnrN2regGUMJoAOY7NFAry/zfKwSlRHxhu
DYyEmfjIB0l2+LbuLuJoY9RjqpgEMcdCtFLbZtsAzyIAR6zKXhDVWPiwRLi/QkgU
hNSltw8sy9B9fiSgN9TvKJ+73EhemdlJrsVQPT2B2OXIAcjQg05DF//JWHDEFyS+
Pr4VyvfpE4cMM6ic2IoELC8ZlyvXiylCMfqVtV988rJ6P/ifiq/qLJHUyJauK+DX
ILZy0U2jPewznyuZB3Ox3KqfRMVbWUi964JKJyqfw8441yjDvcMIFGefJluBZkNn
lpLHKP28Qw75eYgnTm9KG3n1uh3Qi0gioNoSlhXSYQCRMcj9JJkGBqgHMckONeR6
rU/O+NDoiAMpuMkFi5evLgL/rfhYfeq4LlNMQOBH5NCsFmOg+Gt/OkUD4/Hf/OOg
XwHm3lsw2qdENeW6rpC1WSwhOhpqzg0+Ipl8QiLvRHJUwI4jA7HF09k/6AocpXIJ
cA8q/2jBYNeHk3fZQzSHMnFItzPBRQwO3Bk25LVxyPDCoZ2QbIgOjwxrqy4NlQcN
kcvfxmSCKjldhsum5vJSbBquM7h4zc7Tk9WPJlKU/qD8lzC75TLD6P5/gGqpTSce
nKNsu1Em04yhjrCvXGvdeSEoUcfdUyfkRIjjOcvNpBoOxNFqrFUSe8qYjurNeTVT
xR0ZpNsc4tbp8VveHrRQ8X1Nn2A1VQuVtGARxVYyAxeeR1Co/pRfr0P4n/Dq1Pzx
8DXO7MtcnuKorBflQrcsGlADIVyqa4EkRx3+mwnNWKJ6BIg3sfPxNkmFs6+BW2aZ
W/Sm/a+cbzZdRgXd9eueX9wayXUAB8B5FwZ6BRN+ly+qNUEhZbE7hAdOl9Zv49Wp
Yna9UHVcQkXnkhHidIghBrSjg8+Gr55kk1tvW2yP1GfTRhnjUbvIWPiGAc+sD6E6
QiSfb2Nkh9jRp4QHYupUm5645PflLA1W7l7ZlJN93mFSZ1AvnoZhTAMd9wITp2Sr
Qn1YcHfnYDfyZMdC3yOwS9fVckSRiqVZQOmSAgxyL+Fz091j1l46H4lUT6XnTdvd
M3uaMmYuC0DDTfqLbkuLJQ69bkpksuxA1WXSkuB+vU8uiG8EUuu2edlglVQIR3Cf
iHHCxJcipKuPRR4WhJVlCLBaOkT/qs4DDww22P0WCzZoyAv6oDxu+qV+U46HN3eP
qhXaZBGuKbppxSgVfP6GC9Bp0uOOvE6Qxp2YCcp9xKho2bzdR4OcL3AOwej9EMwR
85pwdSKSo3voCo5uAYDnqur4j/70+yq6d345XvXVBYlJaoxGQBIprAXjP3xuStB6
lKiHn71NWA0NySJdj7PPMPP7QFK/45YFfUBqAOC8MdSOnHUw0wcNpq/QJEnyxP5W
ueQIYiu85+s3TZRxH6m9aOS/60C9uAP1M6yaGyRATBmHnAmldAzTortXnOCiOA0H
HJhLFho5ZtZQ0mjmqsJ2prV6Rk5ANS/bvTYlm+ozNRwFQ91iO5fJ3JVKGe+Y5SHc
jZTEFVViLO20GU+kqUqv+zXURv3pEoM2na3n193amsNbSWJSr0tT8JVz+VFZGcL1
xHT66jG9y3cGRhrm+pq6oKrLaLBLsOehC4g8dXFynYtlIaNPQ6FAQWc/PVxU0jUe
YYKjqfv27k8WsFDZ/Y6X2MX3IPZgDV1PIfyk4JL3ybQsDIS5f6D4bK7mAfAPvyze
jbv3+tvzsBOIJipy/bpyZqhsOYsf3V2QaHlTIp+eypvumv4lU3zPxsroiELt5Kx9
T/rIZ9aMhbTc2yJQ3E68kvxP5SaMpCoxkUuo9dxSY6g9JYgN3eA6WXDKtAf0YPu2
cQuKVLIeNuW9wFVLDCgr7qi+7+Px/HqDQ3jClcInXqiUKpdSG9ZF6WQ4Oi8CQAk9
/1xohS9fnYoM4h33OQ5RkhzUux050s4362P2TTo9+V8dzKLBaC/MVRj41iJAEVGV
8cf8p7FmGtRdrOOeg6XgLDe1HjDfRnGwKE/DRjNx6BxZwr8aeRu+1ujWt9xgCFIr
1OGQdPRv3AcvP8sEJVslm06ETu2s5NyHD2xyUZ0KFRscZw0N/6hWt8UTmrOLcYKX
gvRQVF64fYjyqkaYPnsERWpoGBQ3/Cilveqrbf0vSLDTfzE6ojSToj91G4nNAnVv
v2qkS1n1aJCHnnI6fylBLyFRbGYbQBTAMKSaKrxcpN3dOIxWBExeHdwIu7rTJ9Hv
mfbpDWX4EziUCUeE/VtnV5kqpIGulTGkfy2VoJRKBaiq2cCJgpkSzmmU8gIfFFyR
nXKh1ePtq0qeV/yGfHg46k0uYBiHCBvLaoQWQ11fB7ZUeoNIvGrpLPQSm7ZD6qTl
0wyVqXdYo+iVdTJkND1MWUCNzaTkg8+J/5VYzRa/Qd3sL0oTCbq5FxpZCpIUniLj
eIdhnJa27HSLuXkd4Os5MQjwQQuNVsrRYg1QgaGZy1vIcD6TMsZOvAA/+kxh1AvM
XRbPLASTdsJ2bSHyn63eXbY3LXzE8kchbgRpcu70PBKbQ0z/7Ahczzz1IfpP8Dba
UneEA0BeuGHXpMyaObScFwZMrRGM2GRt7E2Gld/N4xCM9A2q99s5MovyTkwjaDBK
UnlGNyZCbGJwWQcuP/gO5lSIFfF5kncozRK0qKoVOGhk9xrIglHQueVv0RScCr59
FrLTj5ht3mqCiBXia5gVS1ICEX1dAerReZSW2FednR8NouAilJRzhkk/Gtl3TbNf
EJyAkvW2Bq/UN+8Q+jJp0oOhjUuE14LEzwKzQvXaFjMTfmz+wYiMzf11CH5lnS0z
Ze+U7e6viTxw8Ax/stGKAUJy20O2Cc9SypbwuIiCbCc=
`pragma protect end_protected
