// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:37:36 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
U08pS7yNh3veK4eYjJimuoGGHLUK4fthZ9Mu4nXJv7j5nbE9hF/KtIFkZaGuSOhi
oxGO3CAN1XdW4gWLG/O3M614Ujys13EIleqyhERPUpWc0/L2RE4UtP26Ow1mX7BK
WjtQoqk9EbDpqekZjavKe1zRbI4GZs22WGrjGaYXMXg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33712)
l2S2kGQValO7UdG7kfDlR+kmAwOQqrKxLS2bAJ1NvpkSgoZK250yG7VsjN9zqeye
mwNUwmWZsWlbx5RBh6eQ+hKaXMznpM+PivodtzuO7OmHg9uDHwtOvI/w3rSUTPiO
53f9GDzGYoxd0/dLd2rnkaoBETVWevnmLxMo19976D8XA9mgANACuRBz/4Tyuwmr
a85ACBYNF4/copFbgSTirpUJQN5I52qvBacUwZnQruJqlq8t6mFurZj5fo04Y0iu
v6BSwr3yJMWNteP2Z1eXQ+U9aVTZ0f8ZhA2ZQlPYBMldiptldtAwqtnNvwJSN4+y
E6Qxusy7NtK0eOWYQyfpl6jMw1efJHi5doeOxbbgGfyM1kD5s9/Wj9VblGNIKVWt
b+6cdNLTt5LQdMgX/KbB5i7X2GBBwuxwKvxxcxgaO4cwPj3Gcg07RFIxhYs/wR8H
VytMqyAwZUWGvlqB8JMwuyrrxeaUrWP8rkjvAthyuRufH84N15EdkIkeKvKKpm/Y
U4RQZWvPF67WZFelzZdhg4yD3bHTPgP8kvkyK8VSuyyobpiPq64NeNQ2JIR3/gTL
gdeXNgJHdsSQ8Bhjk84tPVsTcpCOIpRrQhUkgWPLzltn3EF+Yi5vhJFgq+hnuJDw
fQR/9WguC3TKSLz1i8TatekQDWOJz+CfFrF9KuLCMmRmCTnnDMVqlOmTDKbUqtxZ
9HV+O8XBtcIWuvBfTEvXMus5wK3OjrsePTmSFArKt0o/MpLBrGseeGGYNGtlLvWF
iHRZUOUHz4c7XfM8QUBaEvn5DzXrjETeCOy4Lo5rJU9AKTLuEMi48PClIEBXVJNC
XU2EFA+Moio2bXr+mi2/tmhRCwNnpznb/kIjGzpQErD+m87+FFCPJZ2LcAqG76Lh
4u2SubbaG8V9XGhyqbVRpFbbPwPzevLv8oXvdZ/PKQlbGzUVywbuO5YRd5Lc+4ic
NJ5IlGklKkQh4TPXgi71b0We197Vb3Ya4ArvnUutbxP8R5hCABUzh6s1i8xmRhOS
Yn9Dpfy9AxyLhxK4ovDm7IbWbJHb9c8/OQHVKKNeME9c/y44emXgu9lmNnvGxvRJ
3FVmmhu5T6YhDUlXY8BYZvzSRiyYSqDeCUPMOHA5SdoqHx740qTdQnIwzFslO8wf
xMFBLHU8O7bYJa6S3Tyi4mDwL8sIPH+bEc4vDBO1jZgXFJtTb2OVKPa3g+nUmzzr
Vi+RakVruDtV7CkAT0CVrGyR9x6B1fJDKM7WppP2SwHyw0HVI8qM6jhCrwDrFwXM
8L2qnyIKnaTbJ0K4LldIu8HynTWOtnBAY56RMOmt7iJW3jVUgBhNxDWSRRcr0wPS
bNfLtctgAgk/AwRQak+MoMv8y9EQITd34IEQRgT/a3IEiMbqYVBWRVgaWzzhOh1E
XjeTOZZw3u/YFYsDdkvKezoXukMYbAlqefkmMtv96fQwl1rdt/R3m28akETL1oiv
sjDgSO3J/CnArl4MvppOHYr3Kqf8ukrANPmkaBTRciGLpcFblh42+NTNXmaFMc9l
eX98dAgKMcZdC1zBAjBrt3d3cnb0n6rRc1jm1jGZZCcBnDdxWJVbg2W6ZXxCFPn5
J2A+XtqkyP35UAIfLgnWtUzRhhltPkscQoz8fWUt4b5WeR5abYnOqst/mgUl3ZKz
YbdGgohwf5f4RKPR2TLLbO5GgxzOn0xOevJxMsFKl7ColjXhV0xmRncagr268Usx
AuASidP6G97aKord4oEKB/UevXjSGtAuiRvxtvdBOhCYEFfGM7bu37qPjcaTFFfo
h7LNN3zdGv5CGH94jopOo1mvjFHDReiZo49bZOOgZKkCwMPoDCc/zMcRnCSj+zYT
kGzV1mqeH5ZF3OMUZhfSDB8XqVGQOvh1lfOt2Siw+w7LuYI97CUs+5mJG/Hx42Lv
+19xwNpJuFcYW/yXhTCcoyW0CEK0wjA0ZOVaGl+qPdDIJLet69B0qFldZ3Hs429R
zjp8VU0frVwfhYdvoBq7S3WEjuLs+QpAyzxCiPGeYcg/KnhSQZE0P2/TE9+jOKza
rTSQngnKctoy3zQwXPSkwiBCjARXf6cDxzWPyQ+vNpQAQC6+Y7L9DQoYP65ZbmRs
0EziCFKvL4s9dI1d/chRQ+OBHVPH0lh7jBLk2JwbJn+3rxmuKkzm+72MIGmJAr0g
bbBbOqRDnmRDLKxgA25t/8K6SEyixikWu9o9jYRnL1ZKEJ4sj2Q9FA2tOE+eHvzg
4Wguo189rdgAKA04cSDkOGU9UXx/JPpXWrZsO3jZieM6nRbk/mfmActTqYzZbzvq
mF/crZa/JPHzxRR4JSybId73PR6137uAT31rOhFEyRVTdH/yiHCLEko/em0Rd3OM
XqTqZNN4Oo6RBh8H6gEzwLbsmc9Im9uc7zYcXhfOgkxskEfJR1RXFk7fTpMmSLmD
wn5U4QrtpH0eBfQI58ptMbK1YqTALpIergbDyOPHnw1LXOEZAPe45hm4s5JJDYaU
9Zy5mFVo+Ww03S4I5VFY/wQsKaFWHHOYuVHml+0ah4TzkmGUcP8im6v1XOixeE+R
DxJe2u4fGU0dnE9hhDdhXRNs0G56vM+3wA/tD9IuOt9Jh2zJ6iaYwKD9bun8n4+H
X22hypTANg/CMDx+3dV73ddZhakjfOGLptj4bz0yVIix8pnLxT+o/Ac9RBZ0BrID
DyB+DvxdU7RJfHOkNEc9N09Wp+5TE1q9hJC6t/ie+Zks0Rwt+0uH8ZKx5WFZ+gyp
s9ppYzXH9x+tenBQscJUMTkMpxzcuVuhergx+AZsrocIVXJ//oN157HpfSvGDjL8
S0rtbdECt6A7RmbnWbbED34MSOITXGLlQn36LEoVHnd1VYfuUw+JbIEflnAKcjoO
nUulIwYXTg98U6vzV89lplhy0+8F9LKoVAVKPcZGRaeJzsBX1CuVAb6RlcToW8Z6
0Pfn82kuWOW2sekdBGIGwWGbb/e1d71AnZPYVfVl65yCrNECTgfmHkYk5V9dqqdP
ikzXI7dwgeeBOC5numtbwtr6BLdyPUWeCyO4bWoselgAZFxTpWdyGs0hugCgZ8ss
99GKPPQP4EIqpVz+Qy0AT8wcSSkFw+qTpqgdbRW6ob6sXBBYzErtz1v3BlyjA6Jv
TUZDSzS+h3Yg58guB73hmNrVLoNkYqb576FD4odPSPY5VbhssYZb8Q6gaybVkv5u
cKCb+5Y4eaxLXiHlnlnZDXDR1Kb5o6RLr3jYY9uo/r7SwIRCLpfNMojh75OkvTLh
UEHnuSGyNakG2JJudSZcQPuFt7ghQk5AjE8SdU4SGiXYfti9sPe/1oYGRWvmRgow
bM4N9djH/a2z+m3iE1h2frDYNxD+WA6dILT9pqDXI+YX0gDjUnIw84aqnAJ4qQ37
QHgpXbbrD2b5T5ZnsgXxePq+W3j4LX8KwYnPEIA1fFPdMrcuJH7tABsgTOtc2uY1
m6F0/Qu0Etkms/D9kmHUpNC2NTKui/KPDVOEZQlGosG8eambO9Tu7EY92mgDbR92
l36iqPgp8GaZaxcRMK+UJRQdcZMw5rWvYN88la+pBFLvJNrMx1/m9oJOEy2+d4Cv
zo9zrD/6Q+5r5sfZ8qEzWtMSqbWMgINUIu86HyAtJIDDBD50Fozm+jJHvcx8JQjx
on1Bm3frV3ENQkC2/OQ3WEig9KMofQ0mpD5aTSVMpAefefbgEx9xSLvDSXmWyODB
X++l4eiujOxK5wimqp7Ja+yrzhsn400InekRvALF2Zu5X4Vy2/TCb7YXZPquUr23
zsQoUjHsTc2WvbxkdyX1uDGMd43l4VZUZIA/Yrbdz91oMzhenW2vlsuFhcSaBCgD
/TwtV/4VezjNszQMiQbTK5lahvV9mIVg+0PQd7OWhFz7QUzfU4UzGk7hfTLjho+h
/YlNAWiMaKibogQWXwh1fYyK+mNKnevBRgLe+vDcDYk94A3pdP71+5cWdzyST8tl
wJJI+quW7bMsQrHPcRiVuXZciyXrCwkGq9+1nevbja9o9yANp5vESRlYqCxXIWTY
nex14abVFzinQYXzMLGzs5xu1GhzM7F3mL8dCT74r8EebcMDWIqhEoW3M+i+zxrh
YHMnoLQ7t+XCNGLbQr38gNeMz7/U65e2aimul+kWgF7Ko2ZOvCeiqZ4eLJ1uHCYQ
dRYpwfW7ZqcXVurjcJkvPeev4AL1BwDAZK+3i4Fy2MUllJMrP02iiLYzYGUytu6Z
DXJE409o4rkzVqKfrygQLXItGZsESqhpfElh6zFA90U2sEUlgsphttT6ViX25HQB
vPEUVHpaB5pSJZtLKbq/Zg1+uUoDivUrRgx34RF3j9s3ePxENa15EEJdMQunZyOv
DVK0Fc6peuxGd3hNoM2EoZK2Ea+HAKr2qV0wRWC+wUloQGiKxp10SPW3AolzO6JN
VVwIIFvjKxVzYOzF6BXiTz7ha0DIURVOHTZn5GUaxeeFdGmMK/rE/dKjKIyO7dSf
4nsTnRZJKoDERRb0UjOnTtG0IWA6N3uDZeFu6jMnVqHN0WeuwFH24at3aicUwhr6
ESP045f0mCkrHa2Z1soe0H5ue35To9XquuwK6hOM5gGrzTFZgTBZBiLqCwWn83LB
yUf4EVIuJtcPLjdzWOVf9rWVJYKBvdD+m9tKhDdpis+GD3we3B/jOzLKjJGqzpgM
CCgr51kKeYWl+mEX1ztlCc+3MZGmG9f19fOQYEgZpKiAadwFwuEhciKfEbvkdiXS
tb5Ty5stqg6h8SyAguxLTP7xQCZ4yxPiDs2gL5rsPX302Yg1Aay209s1g+YEK2jy
y2W2XIPgPdc4WPSTCZCFn7dNeTvHf8SHgdPrf9mnP+fNgnKEvD3nAkQ+XLVbFaoM
UHeDo5yl5EMSq+fr12LPqj/28RNrRCMTiBVPSia0Pra9Ubg8lnpQEmO9Zvuza1AF
ooPDJwVyT3uIlcaW/dm1176SyNgO75W6EZLiC6SwqMZgI9pE80txE4qfymJwzXT9
+FjRa3/5xFm4vafzqK//G704BA198tcil5xuG06+6ALUbSxwXfYU9koxS+DUAJSW
dy8wchHAqKlBESC2ZgvrJFRKkGt7WazATQ/g9xFOVcbW005GC2E+LBty4Ozm/hfj
8T7wVJbxw24PxKnzrH/U/skz1HHC+q8n4qO5NTOAQaekWS/nHafb3srdA+ThD9Bi
eem0MbbJF5uWCktOQNpEAsRhkM2deuFPAjQrdl2zJjrV7jRByhChIMxCJtgS6ljc
oEVgcBbM7qgmUezixzbXIeHv/C7dy/gYjCv6herxCe1nsmhmNV+SH3MpNwm9n98I
LjdmvAQm1iVXU5kB3ALwI+0ZL7R0+bNq/NAN5tfWget9I/MiiqUGjqU0LTEla1A+
kXYodEDKDxFJwkBpB7v18ly1YwUPyYetxL7u+dvQQ8EcPn59IExWHeraEoFgGxCW
hJGKBMDKh2qSPqDbflZ3hyKU/8d+6sErDNABrke+b8kyYZ+hWQ7k4f8okxOiUd5K
+nUWRDD9MHdegwCnrRIpccjcwn7CH6DUGuac07QMgWYQBUOZwmk1SMr4KM3qMXfC
uoHFF/aA11R9cnCc8yBTsvb6NO1qfIoyQP0V85qvsZ0niNNLiE+2aE6rYGlrfHuB
gguTTjh+ahJd2/CjLxf51hgzTtux7UAnLTE+SS8X2fDkbhVLO/Rytmcyab2ZUAmR
y/kLgidGD9E1eaoOaVdtmSHSG08j/h2xZDe0SfsXcAvviwEhLM7ldwt5oAgUNZ90
CxeyTFUHGsf2XcTEp6kKMlx6+frnMaES865LMs8HmsSzJLou2DZ74itbdCxm3JTM
7Elvqk5zbBdvFAxqdxBR+ud5E1oTtZ35MBC62EqajtEQHxxu84Adm+TgHUhxatip
gplwHRkLBZmfsNX1RlABjimssuBV3WXbdHOSkhh5syg4EhNoUa9PIGbu0+z0qZ3L
/Pm/xMfoK9jtKxxNOEr3nU0teD7T9IwQQ0IFGL2RK7jf+/9DedoI/LOXvDrPQErt
d7Yy1KxJ6HwGa4oMWeaeEczg4Ry9ujpv9a9+HdwDHA/y8Vo1QB1ZiSRhGwpYicrl
uSI8RpYn9md1uSekDulFgdUVxqbAXoK4t463NzthzdmpjUktH/6MRtDWFSwHnCGu
TbguSr+js61UjdIXKSpwHuciyJ9ApbLc9H9b6m3x6k8xTTB1XnsATnw/5YOz8AHL
FvxcJQ7RaQm3mGaynODUac552j5fgUIgAWvULBK0CPnljdoTqLvAzflNfg7jAhfO
a2EFVUKv3x/so9mAcQMMyio00tLOJrM+eil6FHlEuTeEvsxre78fsJMAG8dJRo2p
S2Onj8V83pmTB31C9Yv/RspJI6NTdKSr8VX5n2xaEwIS+M5snniSyuHcr2PZhGvF
UvifmQPMOu5SGXgFkGwTa1GNJWUJcceil/a7eE3C29n7301Khv/XfQ9Vspj0w+9F
dzbtUAg+YGI+BMI1EmVMwy7qJnwhYqPsKHPlwjyXE8u2iGsHZgVpqx4bDIVU0oDp
b5IQDgyKh1n0vf3T/0WYnbGIjh1HeRfK/+gvj6IeWc9o3pOoHdDXQ6xRUBHv4KbW
8E3HvCjd9xYNd3irgt0qZI9EubDiTd2aoqHVCt/sSwnji3oTHZbNkglnKCGGGNxR
pt0Txk3DHOu22VBfUGwtR4XUxWruRzk+Q/+lkMj9FZiQLcKBU/joQF5d/GWEjP26
X4xrO1NNjMz4Cq4CDhH0PNNwanTgpkN8gtG7oO2SC4wfhNjk2Eb1BXqu2d4hAwt3
vHfpk6/fzcFs/ti+WrxhxD5dl0p6jvjPjRVoPGIpr4o2jdf36Ngrx1GLnbqIOpxE
bXcG1bUVN3wIOoMjzKu8aDjKpSxCeymca+Lttt5ZoNiTB5nHmLaUeXz9jZ5JaS7/
ADa8RtsnF37nucK4A6GO5XvptcNH2kCCvqb67kUgWmYxWjDeQE/pCObYh+CLib/9
De2awPAYQSl1d4F3J2SI4H1f0do9MWbZBG3CmoQ0H3BE5Xko2TSa3WgEtvklZvgn
tmPfJwrmSFFj7c7PW/7jLsktxDcLMHvsXVFTrvFKS1jbXhGbOXP7pi6W7MNIuEJh
Yujv4p96J5ZvouIVAObXkd79tOzIerpW29q3SfHJkTvsfaFPvhEcspdgZYe6WN46
zf7LzUAyDe5ydjaz1u5pKvwInUNfHgznQxASIUg3yPuO65lzxj1Xbcc/jCRDfVzq
W1UygVfdoY8lhR75/3xWEJyFVI/LBrw6upv4Z05p1CcZk36yyFN0ypXevIYy7zlv
Q2y9AI6hDwxov7P+/OCnVM06qEh1dRs7E4/vsknDnbD2Gj1c8DqDCVEIVawwcKOR
tVWs7XdnYdb7NAyX6kouvSZCqZwCL0I6/66vSaUITbjaa3vQdI2pfklnQYPe3cos
nZy6+o6dkcWVz35fs48Wi2xW0OMr8V6D1chRoDxy/pnY1JksN5I1pj+Tjq9O3eow
L6yiMNFZ/HQ47r/cgvxhLI9aLqKP6axAWFX1+dXn96SeA/p1vVv2wQtRI0YTQatV
3BBaZJxV3hRdRnMl+IITAel+8KUMqL1n+mIvitAHq8Fq5/JUYcdcK+SIJQFGJxER
qaU9gHGl0EYG3CXDpLvRt6P8/gUCfjhzdCdEoggOQjzPs9g8Rhd3m2X/D/ZlcEgY
eWeFPhR+LE4Nl4yXql0vo3AhS3GWwKnmXtc0wfHUqcYcVLL9/e2Ocjs2mecf8SvY
uImkhL95oZIciFOJrgC1ce2nHQtiadEs3NS4JMi9gHfEieCC3lvW+l3k9bT3Q24I
dvaU3hAu3jHnqq8y8Rny0qAr4Q8de/v1vgO+ywJrsHZJGE/Jw6aRntFWY8qTDtoZ
V6jUPZ5JA3qH+AR9EwIYwYYrEvNrKnWo0WTtoBLqYTfUeHm7TtidRlyha/gGn/3/
r+OM09hy2GmN1k67RLQZ3z/QfOtbW2Hrz7fJgZ+qCEjIiT5elLnbuRqrOiL2q6N/
5g42wjn+X1LhjkirTBEDJEcGIK8eLXIbHw2OZPWY4aiWz0pk53P2nuvkWgU8k3vC
d4aVWIcG1c0e6a4QGTPT3TP4tw4Aa9LQ2D2ZCY2ZkGPzdUB/T9VH8sUc8tFgnCuz
ZVuuBDRNKx1Trlt1yKSRK9CbbtYhIR0Q/lfzz4EyfPEd3WJ/8rhg9ZEhEYKssG2e
qQztwESNqFP94OU+VCIKY0jvx6QWoPCRT35ix+Iy3y6gcHDJ7LTcMcqc94vpk6ZY
KuSdzcQz24zBpcSFik8eV7+fxOZqk73heDCD1RrIHt2JViIgEx9Zn7RVH1rt+d0d
O+j1q2NJCMFi8lUasjnQ8AP+c+txcZKcia+Lly+OG5wThhhBGxaNhs6rAMfdP609
E+e81ROq0aampfh8Mi0oVHkXXy6kJUfOq81UfHzTS5eV0UhhmB2bWNvjM/cnBiBu
wMUraMSzVFHJMp0jC4D4iRQBOucMKfPO2O3SoL5P9kMwuQo5e1RvR2BcR+9o/BHn
3M99Jy4L1Nmg5mQh02J/8TvJJa6RHbQi90KpwS5LMDvXgi2tdn4GywewQCN9PHPY
O+sit3BDvUA6tSPgiA/jBtRjWB5ZA0uZ+9uBc+BDpbWoMvp1ew4YNVIvXrrOOEXQ
LVgPrQIZwJthJ0twWFFz8bUiqvQpY3+iyftjgQJ84zJRGMCI/d1RJsS+HVjD4Ral
RFLzdImpkssjjVMH5ad694opIyAEgONFUz7XPf9jNOZyXY2S2Mk/v3wVZbvHjVOi
13s4tE20hZBe2q/cB8k+ltlsWQp8xp6yK5UWxMAhql/ZM376kRm20K5/CAhN/l+n
r/7oMu2kBYc707WG/lsQIV2HgAJn+hIC6ZzZ88kgLrj8xRrVcdA145gkExd8CVCo
fQZqXfKzFBZplHydmJ+kjPzJewa/U2MmDPfNVMUzvMcSvBF/ix2ogqX+MUJPwbHn
d96n1lvck6/qXQqERIU3o+ntKB7REicbIVxcZPcr+4u6KuQTNul2J09NeCyCWP5+
DIxi+0/ekbbwQFKaIsKjdxakOpIMIwDTLqaIXxlVQr6paX0qWTWCaOAPnesAUCRO
7+BRIV5A6EqJ2QkF4kKet9e9JXw2fof+QOse2Wi4c/FuIxpJcFkoXvExGHL/vpTl
MyVsoY2TuhPsLKM1eZn8lLISq8vGlrHCOYMiwA3iigykeepC+fOXU7vyeItV/vWv
ryPc6KrZciV5g08xopea8VReBJ3F9HDLYXABgBMbT/LdKFfdARQo/JAaS2smyAwv
YpdvZlnYH6CrBn9RLpYUz+Cz2wj+ULxBvSse7dvrB+ytQVfsuEfIZ5qPUqEnQ4OE
BRrNUjdGLNZdJgkubNUD1QJUi4tB3HrN9v2G9oPj42L9naxGh4bYSOCwxoPvdxma
tiYKgnpJV8cHECmIlNx+eUGTEcuprIy8Z/NSCAGp9qloiCjMH0TI6Ftljr2KzSd1
O4bU5noiDL9TEPFNPoBBW51z6ar+BttMRMCkXxNHBqSA6Pi+XabMUyBlS/oIibJy
uIp0GJftKNVHhyEAbpyfsWGkTRdpFG1d4oPNLPdUSfyoUqbeP7fOfULm95tb44G4
YqAS6vDkgQ5i7fpggzX91FHHCe10UGcHAK02a28AKxrNFkiCWPdXjxK9o0tJ5WMu
SRr6DKLhDDU5JXn8RERgdMupeF57Qb0tk9pnnFK1Auv3OK00vua8juhV8UDNLfX1
UaE1hay/KlYu/uD7yk9yQp2ICbWOzDvk81r2k4LoRYKejHL1L/lPnqq6pjAX3ca4
OonjPowHHlooJod4v84ICuZ4qhqAg2DH8iF4ATo1eH+FGmPWkU/HFgnsizCdXrTB
DWsBPf+ro0CAmpYYPDlPxqVvSZqINg+awrKxe2ZNohXnIT4P9gWZVPPxyZRBC+nu
g5k5KPQkH5Rq5Mf1fpWODInQ9xyt0Co3/JXaoYjSoB06klhVLC3+KUynOADHtAS8
sri2FJYmZFS+Yx30wQluuVMBUK6MMvA1SOsJqzy1KL3YuTptDiDDX1ffleSps6py
nU5Jq6XmG0sTC3E1JDMhVKEwhrHBkwv6G2aElC8E6l0I4fb8Nxa6x1Mewb9GwyXe
Wbi19cw468IOmT2Y4z17yuXiuT5QKghGQvdLxlTkuKj3BT21CnTM8rijuzFTyKFk
XLqkY0fxiBIRJ5JCvf9J08GHbEE1pjW1BTVIHKoVe/ZZcPnj/UXq4dH8AqMEv+8+
NC5EKzfNULlyFVPAvT650AOd7oksUm2o1Q5iS6SFhMp/gTU2In8gx+OF5R5xS8KT
RpH9aOkt4t5Ce0dDYV6wq3385MyJhXCN8lgcogdPSwarXDOYk/AjQHqtDBvBcgrF
FKTpQIAp6az4dYQUGzorNEeplGeZ4Y8FjTxgZiTkiU4PD/n74N/6isujqIqw6M/U
URG31j/jEDfVbTMIWhNOVT4JVhl7eq9B7UixJ2XkTmGHqXBzPQhFXdFGMUfGnn+r
U0+jiq4BBGzucZy3VnQeUYoMzPXX7uMHjdoR/eT7EvFAqf8X0i7Wv8cYifk6kw0/
1HmUsx1/8GmllTa4ECwBgzHxcwC19HfI0KdtroJZcaW7s/Uq4LetB1FIvKlPBXMT
aoKcRqdLdWAvGnBGZueefPrg2JxzRfwo1u4KxzzgaJFEUSZ9H8PRh6a2ev8Rkw3B
prRKMQfKSlv827mbi/4uzgTI3tlqyk9CE9IwEQw5pjPjGKakW+0f7Gei6JS8ZaKb
wn5sMvy+BAvYwR9xYtJwyL8ubStWg4hsa+z3Ui/SbP32It5wdIgHOUaMwcwQuOYm
UD+kguGgmIQet/4+TRpDLaJMhKx+AW25dpfhAGxRPu5kpyePtkLahZuusXqsHefN
gCGUWbt6/qUj3yI0GlFpE3kdzMyvFKg0Fhaf/bGw+y4Nhg6IqLKGKBZIFeML5EYM
jYWkQHkLNtNHVGwiNT2aRz9nxAqXLIrgzqhJ/HU6s3Z3YvfbTgzDdsvBG6FzufmE
5Wb1GUEFaozQSxDi+kmaimZFW9463ielwPHmhRXV7dh4IFX1NgEuVpQILQwUN977
uMbHbxN1QpEfv2b+pZmFKEvMzg98TZ0kHuoIiUVygRGO6hpDIPaGfgAcKWNMifwG
dVctJARIGDD7faNtVy7n7fA17CnQO833qfrNtLXtgZFPXZzMVt0m8ycxc+HUqBhy
Hbb8Uit+ehR+iJiHT0DlxB4ThXhWyOmP1arIgXFWl2N3TWW+WHiNNfBrwucNuxbt
1zsmH3ncqC2LbNvgURjj1pSoZ4AhDHVBNoqHyeUep40B4eTyu9grncHmeGI226LI
KgAqokmcBwAc/gR3xa+3NdpAUq0DMu0t2BipzQpseLb+9gN41BwC9gTqNE4WLhmK
zzK2TgywuEtJNVEEugL9S8e/LavfZFTdYuQwbFJz84TL+lzUvuI71JAMcrQ0V7OE
UABlvAsZm3hI9BRUajjKW195rs9KFYHsfC50oAkcRa+JE9LC+lbfslghTgtwxDSN
SSZhKwZ6u1wFi80ur8gpFcn6w/Hj/VZ0G6TcTn1JcP80udNfb3XU+dB0tgfQxK7c
NFJkSCTCASjxYo3lUOOfk/I53ByQtkWqtGM+x8JyA91R8dQO0Zxt2O2TiUVOKaQx
hsGqLRjyFOM4pssqP2oxaKdKHnRJV9FC64pQeI91u49Ldz0vmOJqJV1anI2mKykd
0LAZzjEcRZHLqirFRSk57z/NFScCq7kzxN+9ilyAM539KBOguYr9+GRdGNyk8+4A
iTvKBOKtpkr9lRp+lrqbwViTkJt16epChbWhS5E63H8/aPQCNG9wtpJPo/32Hw9Q
ksF2DJ2/kdtETGQLpfHjp3pbEgituwok86rgsb+iaBqZcYvzM/hgVvkYPOke9HJg
MbkXqwTLxRmiItJ47OMuM8QSfvI0HcJQh153TvATKhTWcnORqGNTXnqe8JS2P1FI
6qnKE84xkTVJNjz4ovMJQRdmDqIUXA/seBxr2dPRJeXloosEJBrBXwgOibzpbU1m
7YeBN8R2n6YE47vhiYHElronuHPR6j0ah1pk53JbEvxIOYH5P0+uUv5OlDX8xw7c
71WfteHBiNxzhUtUV/RJmg/9+5b4sxXxM31V+NOnfEmcplI8Lq7Hm804ct0E9UNT
KAX1hcWQf6fFRn3KaDj6EuMQXX2iezNWaaRZzB2vNJRX/uljnifq5fUOrxH4Xwo4
vZme1mcujsh/fWpuIn8QFGn1JyADCOppvTC9P65f0Ut/sK7tMqtfXNhrwmduHU79
8DepnLFm6LApjVExwi5C2dBSlcfaHlAdaI2D61rTTinuw2N9P5k4mpJQHQIftvFy
9uXYzI1mh0MXsAH6Ehm8lIhkWaHNQhtCWoZ85SOIEwjaIr5BdKM7yyOZ6qJTQegM
bX1U7TSuTNr8Xmdg7Ff9FpiLyzUx52h0nFwQmlqcdkftGthjql+ysK+IFQS1K4HW
zxZABtFYSE0YC28D3zKshDgs+5ZlI2A+VW6i4rsUkg4WOfHY67ZtnMeM4uSZ1fqF
tKsu6VtDfkfpNZC0xCKPhtTGMPhVe95ETxkSaqyFkboHLgCncqSaGmsbxhqZl0xR
+Xjm7vnrhr3N3kmDgBlFh8DmiK+IvS/YRFvwycLC1eU0egb3O9gCf+wn8XmJhwIb
Q73f8bVGQOZksRzT1a1by65Cq0wbaD5g27lpycjDPIpVy/RgcjeVc9ZW6+CCMUn4
u8ZF2R0qpCEPzILMGdPQR1PdinYJw+l5NfO0MfRHDxkVZvdDfMZRBjqX+O5erH3I
KAExswM3HF+U0JDdUejFBqcx9sIk8dNLiGvDfdgGMR4+1wQbtuzJpEcGc5Lgi6YA
oXduLRnwJiuBfqsZ1Z+1WJoZV/7B2Qte40QRU9C/SJswvA9YFdY0yYRAuuWwZCme
ex5ugcdRY/SmLLIMDDkxojyKmA9NEWcjy1A9Ab28ZnrNtHOMT7BgJFwYS4cARBxm
8YCbiMPN3VpPCkia2KenOt+5K4e1SXOQunbbDOH+EInCPJOkdRjykavsOimDzJIm
bOtz5X9PwJpZmjyEt6f65WTV6VglrJa3KObYQ3mRKSrXks/0bDx4UMQW/2jhY7st
bhkvBz5N9esPPiOUaRlkXzGKlyKnj0sTHUG9KG0DfACvxzFSfZU5Y/R+Oz2PwuRx
ElO38ITi3SpMnmupMpCrNXtQsulEPkIZZN1yBp1PtescnFBxdhQzRExWh4PjChH1
uqqLnM6xBki1D5sgopB6fwdCtTNeR8kTy8MMsDwHH5/qToWvudmoHMFO1X6xqCCr
CEj5rtNQ9mGeZVhOOWL0zpG7EZOadzCT1kur+NpebWBy561tYRVfJZvQNMmgM2e2
X9AbW7Xxw5ZYhFbDQdWqvw3e+uwqSl4ltCZ+UHMrF+YbkAQUdb7xxJ7wX6Vm85a2
6CbBHldxCKHD9WXuLoFeW8+1wF19WQ0blbVESklX4CyEowvhHegq1j3q4Av8fnRw
4lGqbFa63xSW09JZ4AYTQJrsyZLJoxXZrYbAuuj6+KR26JlBB8SAhVNnRomF+El9
22r/9NdU5URlfz5eOoaIFdRtOOsNNNf2BeNBfVuFpNlMsQ0XEdeM1iIzG/+zDZ5V
b4WlR55VXAfLyxAuQ6TmF7kM/hsjR0kG0wqKuf1EJaAxuAK8l1OCBPR9Ypi83JC5
bOi9qz5DC3sMRuDELP3QeasTQnvF6HdIBK019slU2nkLzSEXTaAauWtEL+/BI/wY
RIzSK/AYbbDooodqBsUyE+us/nXc+jU3A3lbn4TV4FMLABaGR5IKEBQDbtPFQw5t
9cSsyKokzZlPcMYXNaD67QMWQFEUanBOvXptpHKxEb65QbiyMpEqFdfH9D/HpSmb
mvveIETn2Ruc6TgBBI8kTynFfZ+BOc+rV8maC2PK+3//YxpYZieiKPMAy60AoF5B
8VuRBj81tB1hZ+LtGzcAqT8/0OOKAop3SWNMMDmtavHZ6MAa/NfglaXkddd9OMf1
YobVam8bZJE7fw2ksFPA1ylnhO505z7pJhKamthgd6AOovG7o0zSOPWXopKe8Q6H
ASQcD5t9V2oO5QHk8gkWoGzYg4l+JhEoCjCmDAyjZZxOfQwajfrmw0GzwkeqklS7
fL/wtTj2miBpTUnuetS97hgJ+F06Y6VxCQKrj+8M101F6ILBuQFATa7LMqbj08cA
0nAUbEWXT8EAIkg2P8fPWQci1jtWT5l0pPykFPfg0rTi/vnJTGxZ5MxVrR4L5Z6b
bG2nttF10NGeNMOEOYChgZI18H2OJr+XGhi3PAcuLOIxyKHnveDImg2613zC7TR/
AsC29M70Mmxj9F25L4SOjXbsNZlnfm3KC/pZzyW12iMyzV75TOjT01BRBZnRKsI1
YRz/X1+n0X85uX0VN4Jnj3eSeQ9t4PMz8DoUAH0jN8GO1QIld79vy1iRjUJYY66f
xFhz+qtoLWxIqPHxOt96M7SqySQwb9g53tDkb8cVF40iiBSD2G78NLQgtMk/p9x/
5evgimN06aweUMSJJK6jlRL8dYpOL6HXBeLDOImyXNA1vbz7q+d7Ks7JNvN9CkBy
rydz83bMnzOozTwb+WjAiXGf7lLavLdnfgfeqLImVIlf5bP1YhkL2tztLiaad15T
A/v3UA7dCmjv8jU+vF3sJVjYaFsRLQN/dakf4DtIH9TyTFMnVYkMI6UnZ9V5NJKv
wtAg8c0ASmKyl2inN98mMdCYg6tEKtkossFKh062EvVJkKJ0ot+k4JqaA1lOGgvf
M9fJN4WSqx8GIMddy6k3ma7akUTG4sMbhRuin3Iq/MENvorQ6wp1BOdAA5VwKxdD
TMRLBexkYc8jJi0eoVteHXpQj2gpm8P7Fm6MIhkHUSwoT07YrE03ij3+MnlHjvAP
WnGsMBVS7aaYxloLNjJSY+Evbe5kjBjS/YIyVw8wiwZFCQjIfwCPUeeCOFg9m7ia
0su/GJKgy18KjxhPsoZa70DrdQ4qealRA5q0IeHoWlPTRZZbSS5/VYu+ZQDQrLl6
5qgPbOAQl9eWv57J0mXfR4NwR+ZP1ikr7cSZu4CfZSxjpE3edmESRoolt6FMH5RU
z6BSZMUmdzCS2ovIeG26fx4jx3ATkPCwY5S3upUQHHbXdrwP4t889cE3hBNvOUyV
IHTPfUMTKkd0wESAgxchkbo4RTZWhKC+WiECxiukKoJkQis9pOoERbcUe1lHPbkA
Gst0+riSYgEZJ8DOXC8jwDmPZhFAULXGPQRc9uerksZPVRnVdbNgcmxRd4BhVpba
vL9jA6a8bctsLMoxzprVzGKbKxyEOwJ1J15FDy/c/swUqzIkksTAse4v4DYYDQYH
GBI9RRZZO1Klu7L5y9cvnbjfJFyMGRikHJ9CDHRVptFsR2iHXVHz82z3Le6KcYT+
5Z5iNPdcHv9KygsoE65WJ5j/CiQwaG1qKlVuUfW8CcrlacpqgmZKzeq0fVvq3l3I
zyDZJdK6/ILf/aIQ9HfsPdK7iQC8GQEMSgo5ZnOr5LluzUNL/uXZgMHpnochgOUI
GB0cz+yWwvf1C/6Adya/WfdvuIzWmAaW9MCmG2Uyp91DHHRZKZ3tVIouSD7mSE/I
tezY8KgbzrdZSMjkNI7jtei2QcB8b6oi6DUSvAca4jfzjjV/4UBSqYq/MreC5qIY
2bAuhXHholIdchsDyBR7N9wFu30ndJZKfmkw0yVzcSA6gSO7yJVqKmMYDR78TzCM
XcduL3fhFhrucQeVUFLFpuxVCnlpWqve9iJMRFWteHaiu3VnU3fvFZhEtX2az/NT
L30s6SOdAPAaDULuu+hVGtSAP3H0Hy8hWtJBbRGk6ffTEmRXYukhKFq+QCwPwd3u
VBdpWEDuC51xDYFMDJugjBFdKk6G7RPWLsiocUrfjO4tWptdjTadR2r41hKDv/jt
+mwVbVThollXMRx+Agozrgcj1xBufEo8fPiwQcsmvHohsXOyZrY6d4H8GhAtkkOI
/5KZKgObGEfmzh94561WO/QQ8KcX26jCXQ00QAx4GZqdn1QqHnjxC3+2ykTDDC7n
/olOJgSYPk8c/sSaZJRSypV4USE0x0lE2dPux3wsfExE5M2Xall3LGFPEONr36/K
QPvAWwDpEGyobZP3eyYXXDOs085V06yCBTFeOY8d/2PdZRetrm/Hi8lrBIelwtX0
wxzAaRXzf76b+ndY+LiYbBCD0skKYyJaWRw0yrNoJZ1OjHVDl/+eE2NaaFD+T1A7
J/04v8F5YRlsglQ6RttA5Aiz3e3jnvSEKf0+2+WJda9CR5vTBey/8NSAwZJXAouF
VJVQiAHrs+0GeWIBboEo8pRQtFlGJn191kcjINNg0n/cXigw+7VNxIUNcS6XT0HI
Aj89OuNl9wNaAGEJEVIZoM+a1dzTBbMB1/7tdPBvHqJl04gFUaYtHck26AXZohpa
xIKSH2w4KVa3mgxur/psoYJvHbbv92qipy2i7rhtmS6+Qtc+zqfulsO7upNHHDfC
wmd3Hy6cGQuOkalQW5fg1qiLy4sgrJFvzZKFrMQGkGZbCH2THYHVQ0VxL4AvzT9L
umxJ+AZa73Wj51XrO5IJ9EkFjWuE4SBpbhnWWMfZWpIo+0GGQWpxgukKU/F0rpJO
waD7txubgLRjA6FRCdy1BdYZ7zuFd+pu8iHIyKmPLaztj7m8BY6fW+Uoyvtbu6gu
wJPcBH91sxYtrIJW/Uh/YpHgYKHPDo+Exruto+9KCkx4cru5mFtf69K6np/OY2/Y
xEwqKq9YDdXPM/rEWPcINR/ous7Rfjnmrmf0YkW3rzp9oE8zlFcIYJLu/NBVrA22
j3ZpIKSfoEcbqr9Ln/JJT7+2cWpOi8Sehi3F891vlCXQrksjuOjiCkLPJzfMSHVL
ShauTEJb1c8W14jE0HGwvlFb/CImEnXhyLYVMMjAk5actuJFZOzseqZCwD1/3IlA
KfFOO2j9jRT+dLKnfRv8sOe4iVLxUiWvyT0TXxwfrzWpmbGUBfGjZnuTRlodDhnr
4vO2/kt1QHqlUpFB9qeIvM9lP04eVo/JNdIF8UlmMAeDdPuUGpHvefLm4mPDm+29
lXE0GSnMiGqp4Y5vMxkcXqN5wOb5oXe5eKHXCwwbvPSUxkyH2WvF4/QaW7bpqgPQ
Lht7qbwlozQ6mHt7IfK6peH2xOdiALweVgpahN/ebpWBXxqNmv3KWfxTmXA7PjCt
9E0DmM3dptcYgK4/kwLQhn5uS4TbgyZZlETdmehq9eg/akvWZgjrxlX0VIa/iomS
2BUFgkE1Qi3ZxzYn1CoEgjpE9mruvp+ZVHjcuQ1nFxLO6BwlB9lyQ3j5jMiUIBnW
2tyNxKrZ7GQkI9HoPtxjxnDTRfaxocm/006CglnHwMPSlhGWoISuDIQh4HebWx2a
PY5lkcC2qqf6KqysWvsZM9I+tPTLuS1zjfAvi9ym0hmyQCDKofQD2ZdaLuP4vJeW
zNWbDxnlmEmt72t3w+ACFH9aI0Drr6M8fSrK4lYAsOB1kHaaz3V0+U0jIwgK+lzk
4FLDnZbqVmd9o6IVAcSAPFaYXkBDI0vrTfgaCa9qcJ2cTYsIMjQ2s6Z/U4HfBAW5
yPAD5dEKAIuJ+zT/cABqjZHL1ZW/ZBGjcO93h9e4mb1LGDVLw631DWHQVRcifyDH
g8b938MKJVnbSOBOEvvr98f0Q78/7vNA+6mhWqdd4DlAo0SMOTypkXCbDihpmtgb
yjfiKPS50d2vD93Ic5gUckUs5jIX1l6v9zwCR1+EychiDS32/DNfvVMV0attInTS
QIzZwv+1ojg39n8mLgq75Uu0VauKH0nXkhsi6iINktf8wbKJzl8116NEaL4Xag0A
8xXsVBE6DPQwX1c8cc6BGHq3YL3L92O/IhCD3siEFgKfuIwTxQ3aKVl/P37/bhXW
fe7b8eRdcOGkgWKIFcTcdbQe6Ky6CSaKkVXYZM/o/YZ9LZlOGjzl4niS/J1y1jH1
U7YnZCBsY/LO3njFEE/gmnBOeEIKQPHRrfXBEaK1F/j6515W+XxkndmEl8f1cYrb
M6EUYDAa1dEVXesaipbkytip8DcEDLCaoTAAF6posMTGHOxQWxddmW7ZffmOfPf/
63j2Tzfm+DJB2JGrvYJaJJZaN6Uc+mzRYSZf3QeAe/i2PE1z/N9CuDUUIjUTzjFK
dHsaEtLoKC2xNrTDNX64+3kFzQSEDUp41qoNJDCTjs+9SOMqu02LNBfPUc2MeHOc
sVj1xfwh/uLrreWWOXH+lpbAGpCrfMBM+KT19HofHRlUnv8pBhGP+70jlkuEK5/P
mkQvGfMb7OqSz1XGoXi7I8CokTycYwNsiix72cbx0Lgn+XzKi4puFfpF/UWA0KjO
BAZj/XfgPttpQKbHOPmcaS/P0h859pF2FZpexeMYgzTEm8CJToqtjzTPxTf6r8t8
VXkyM+qMJ/vLI6/y+WEvVhIL7RMzJRrgnL+HaGg8R8eJteQ8IqTdfHMQUekHrJF2
EKfPr609ZuJaXRLP9mD1QJNaj6oWfyKcrB0HueP3NDLId2S17dPVnaDI2LKkcRuZ
4L9RoHUL3ApfMF2HaIxbBwORgko6U7TTjZVGPRTnsrsW/DS+u0Zk+bk6/h+7kWc7
skO1RJO+sjXnOn5cF1DBJXLyPZ8SoDgsQu9xDBLQfVMRJPpzwK1+j5vllKLaKy9U
5Qhrcd9xan5R5WhcvRq2XndNtrAZnPhy0ZmfNKVxrlOr2l2GgNfh/bzbXh7u0EPk
yD6xqHaBXCLL8mNFM1/KpjQADdy6IkvurJfrt67dvGCRMlBjcIkTaIv0Uy/7k3dF
IH99tG5FEBDdYttxTzq2tSihrizN9Fg++kVvvXuRI0A5w01wW/NUzMuapY+nAKfq
k8MPSdolN7Vn4if/YwJHKrL/mdHAHOTuUKtWVY0MByRmsJWuq2R3THrolITdul8W
ag9Wiz9nZLN4mIu+FjHkGCLNEiOY2TAEwIm1vLmsn7+ynLcCG85ciJZyRR6OzdRh
ZzUBA0T6owW1Lm04nJV91tfrbm1uxjByn8ROd1xdanGTYMEO9BBVuvBdNU3fK+Qw
nAGtJ4rjag1H8zmi2PdpYPtKMqBbwZUmQFKzbicOM7NwJsTrz0v+ExcXp1lzY31T
U/JQ0kpJX2nEU+7lx0Zfy0A9GRq1ROqwRffatHGZecv7MHsQQUvdhiDfxYAVsEDu
R/iqZYv9uXhxAHZ9Y6QEiNu9pn1EfmOJhJ+6c1ZDIw1AHbivewWj1NgrUsS+jpmQ
oMGos+oqlRVQ9V9BhQV3DFj5EeeilGobkA/0aPtJs2vJTzydG53YjzHie5I3+Wsh
3OAngbRFy2el7bo8Lnke6FKVarMgPqp+/1gnS/Xb60Ph2GiuxzwUubof53UHovb5
5dDFSWfjpxMrCI6bob5wZyz0dgR4gqlL2fiTmIgFzpLV5qDPBuafd7wiSj3dswFQ
NQLuN96F3j9QYOM6fy4Lx3jcCSzGWzdtTnV8Vujc2qK5rzYMGbuHHuf3DnnDDJYa
4VlHBYP1N2Jc0iT6xl7uhWJYn/6s+oKkDp352pYyHiuXOc/WbA/HgbiyeO3jbgCm
MVur/btgWPmYIEgM3tZ6f4UyxlS6fi36mwEeHNv7Y1+tG6eoGNKL/aeDWp4X6N+q
H19O2/spZRIwfTsNWZvOgReYLzXtB+fzwUxbPBqz7gk9uchLco8RNNSr11ti0JFZ
c3BFeRWgxx4PVzruafKtiQAWyR0nyrG8JaVuNyl24JD2W2lPxDzkT6VPqjc65pOL
38eRJhuMcg6dMLHgXIj2S/mKKYd9Ao0HR4SKM/QNyV6E3RcZJI/hU+B4ble0jT0N
XLD9Ps6y91RzJIPskzPBkp/76oQq0KxqZOJbOObzLI6rcyz0ez5TNw2e8qUujlIE
DO1o3WqIoGYQMA2h8Qbys9na2y4el8cybcVnYYCB8TFKPpdBJSrbfsItsdiS+npf
Y5+oIoUJ3QCjDmsro1Bq+KI9C1xgWK1B2fcvBu1Zai9dZIyY+j2hY4wVXcPVIX59
w5c7n7pWC1N/3R0NDhkMdT/iLDtrWnZpsrS2cQGiq5NKBDqcFp6EOHW6IicZpkUW
7msqh9+pZ9W3U4Z2LcvwXG+K1f8lTpP094R+agHFle2Q7222sIgmDI7XQlYJD2Ta
IJg/wpFd9gDJAuYL18QsTG63IH0HmEQ+RREzMsB+FDj/xyuioBAuHtmT8c0g2oGs
/Y7OCGYwSLOw7rkqfaWWCaiS6mTQvTDR11v4UC9z/q1nBoHBcr9wt55z3g090oc0
m7uwNi+j3EHUiJrm/+HJrQBXtZd+pkSyfQTWQW0wrnFiiK/4FPxhPmgY99HNFO28
PglZ+hWpFnG3Mr+EqAINl2N8rauKoQ18bQXIy6QXPnRJ90kvrI3igsYyrvep5onN
HJbbIP+2x9PaBnmkU99uvfJ01EA6nNhicTE2wUiV5EMZ/WU99eXxiwSMIgfhL57e
IS0x3CdyaJtovCxu5aSaTTU3Hei4rtm+qsmysZsTBcxcTqxlJ4DEZcRC4MlY/7qu
cniFu3WMgneYqulmC7BuBF0ZK57IM727wTDJjdW2x2HW6Ed0dwUu/UQK6V7oilN5
lM6pPH4kk6D44cN0VKrKBhjfBrEzFMomawCpKHNTS+LuMtr2A8RkFIzby1VyB+Z0
ZBEYQqS4XYduqhauWy0/aBAFrD3IUOy0b+LzqUOtA0xix62Fu6VQ8IK2tAoLdPuh
AkDb31sZc067vyBWc5GVLmVLnM/AasL9smX1jNeO1n3NcPAHN2l0W5f8nLHZcgQF
D6uuNrf3zQSavcIPCFHd1Ca8ZfVAKZpErVe7dmWXdZ6k+wv5ncloqUjP2SWdWeLc
6o3OG9HitOtEutmnDdHIGywUr5yAM+n0nEwiHtjUiFbVwRAZFiM5oawjw4MX6Phn
EICTje+pllaa4ndGdkdpfWq7/v/fkvM34WrbTvw/LG2kEbEVLuetTGHpZv7RvS0X
GONnOm20+ma6WWBBYp75PJWul1Ad8NC6TBk0AFmdZzWIaS/WYbG9HlSt7hB0jCnY
Uo4KdyLzOhpJChQAf8Iy6omHu4lhtk9pP79uwMbdA4f4uftVTJSUcEG2tkQm9AEe
Jbri93QosIUmDbbwLseGeOdTSrsjM2BqFhACbnbCs+Xe2+EKYvLVyABxxBCGgx5f
IsPfgKdsh8gwbD2w8aEPPsxJvAOzPZFIAL0b603UHljg3/peOpPnBhjSfxbKJ2Ap
7aa7o2/2H/EI88Tdxc+LIteTC2USAHSRVJYNWYPj5nM0qapsBNPZTmN3TMahSauW
yadJnbuUG8dNV7EcUh2KwAKpeRE4yAxzZvmeajQ4BfUC4O3coq3cC7EZ6ZfEYu4z
nHxKCS5s6yuite1zBkoDDn6iLu7Fh6+2QJ1hR030uabztqbKpx9+CJWLFS3oVDVW
FSyBPYGwp9pbuknkox9VcgO9rLorI8z8D/ipbodvd4PVpqaiz0JDRTitu819iFm/
x49I1X6jsVEgz/zn5TkpJVCApa566+k+f4PTcqt26BlxXTa4DsNDdjufOnscCBJE
HEsOxZU0sdJMNavGW7Z9OyLNucQsiR9x9DayHFt1dnExD6GG9iFFcwtBjQxOU14W
mQpnsRCsTY4wVnhbqxQGx1V2Q8my14Mg54TPPJMEBoj1ss+dCkB66BDKF9D0Eltw
UqHPXq5/mcpDbnf+35tMf182/tGYZSzN/8z8MJ1L3y0lgC2WS4QC/4TsziDtNv7r
6BpUdlqhgQQA79OvTMdhxfy7eqdhcg1zAM7UyKNvUcyYgHwJCY+UuzGCCxnz2MYe
QuiR9mT9Mdm6pTcEGG/xHZLihKw4tk4FzpxN70X6BKTapv1O5PwXxXOqunoHdYm0
sgoA/aVqYa/y7rMjPyRFmKa75wLifrcbhHiuL7JOF64OrolFTgYJ9+5U1EA97eh7
tRLAROmW3yP4HmLseqEcxD0krC2TJck43oZxF+R5iSzsVa3AWog+h6s1zJjK0pP1
TpWmD51XdSoYkBUk3502swdVoHEzNgZ4W8s9u8Skd71MQAdXLBSUKrN0K9IJ5k2B
4kNx/1VSGKf6u8Sit9tdlsb/NYnuMF1TXgnWY/fpNT8XK5zKlAgzUTgXWfJr9BLx
FHvkz3OT8ewMpJYGWUFq1mQOY0m3TNj/zurJJoIgojTnCrsEfoAdaPNHF7TsVcEd
t4qnIdUq4cwPb673YzxMs0nl2EtesdLnBt9QEsp9DFZRgLZYqL9ufmQskp2VKQMW
O2YfG78/WuWeVfpA5Gv8CTmVW+NCU97VD+n/6C7gKUBegeCCWaFC1vue8sfh5wbE
7YX+e3j+7dekUqD0AmLuxKa/yIoFd7i8mbABOjOQB8vtIALlFm5uV/UtRKLCy4QP
iu7+6okyjNAN1d/NvNnzjtSgKZxfOeHbh7UxXY0Us1UkaNDCYQQHDk/oH6GCsvA0
Vho8WDMw0XZ2YMcULyZ4VII4ELwEHgSO9S94pZbt2HsTzzujVFRjetNups5uFcSr
f8Cp3afdib2ylJush0/kyPOm5KLFR1cKoaqj6PxpcgZEC/YsVXqoUQZ0YbejUEzk
YjSBsWcLHOc9nfczDUQr4W9n2XHPWs4F8LG1DL6rB/rhDKBOMAk6gO8LrVMe0eqX
z96At1Dn6PlZjBzNRjWVwOt4MiMhCLqwDJtNxpBdehL3glm/WN/jRidyHwpbPjOp
F3OWTpGtfZoEYYkRZxghQOg2UAaHtuXQHxnjRSGAqR6aQ89IjWGmWgwVuZ5GxApm
l8OcLla31N7KpiS3x0dcSPH0dpcQ/klcVKD6Q4za7BCGEbgQMQ6w7Ltsv/W43sYj
VdLGwzB6aYl1bMGDL1VcTcG/nX2aQP6igluw3DLtdrn4ADR11neakViNUT2YrIHP
C7BftFv/k9ymsJuznW12tVopuYix2ZhKxw8Pn0FfcpQRcGVItysy/fYhxEZfEPZu
XoDJOI3jz1rgn74TV1Zd71NZNPLLMtIsHC4HGsj5f+DtWh57vddAgVL3/8J/HMWP
Lug4KpIz5vumSmFcxiRAgNbDbL3EzLY//Wsmey7LD9EBcxsv5BcacgzSQ5uZhV5Z
AODaSk5wJ7p83YXMb2tMHST1sShRgKURuL707ny9AOC01j7cXP6pzi0B4YGjTT8k
T7IxiydEiHdmhNCp4p+GFRoNhLEwOP0CPldiysbFyE49OkugLQWjnD+CkrYMmHkf
nKrGbMbxbRJzlSLWZhSRIXwsHUTAcKusbstO81pX32PBNA8nuPoaeKyfNwHaPu26
RnZX6T23xk0g7PDVc94SnkCVw/nsvfgQcmoDjwdwx0aDbi4yEujMs6Rh0e383HaU
4jUqdWOV9g7irgxaGG7aGiSrQJSCUQ/MW1ePDPfQKizqxJiDRlf1SBuerIQ8PS1q
ZvI6UcqOv6Wd4qrjkXvaY2KmKF2vUCHkU6mfaAl98bWXX/3GmHcqZxjLeMCe7RGI
uddYi8fwu2BBzDV46WBXk6ElNrEEENob/aOD73mL0l/upegelPg1TFHrtnOW2hvs
k06I8uXPS/YKJlm9jas5JskNsrtIDCVhKXM9z2VkmSwYMOz1px2q+yaRNGaS0Znr
PciMI1dIxPDacLidB/9PzHibUfW/w7MQj7gyl1ZiIT5n0Pzolsx9Y/GwuXMdTM4a
dNYPcXp/568FECgkkPVA9wm2kC54qC/MCtfi4dJhXwwJGd2qaO3r20IqoHALa/Qy
wASCnj9eHAYf0fa4JhOdB6KhNpuSwGKSAHrofH0kVvJFX9Ct8vrd47l5GJF2nrNA
OGf5fyJzxmYlzJUtNDqw5ybql4hV+mHMJkh6vHOBvhEfGJLEgt+E+oYdlO3kQ1GX
1VdqbKscSNEwaL0B/3NCZjSd2rL0O297hTFLXIAIuxDcP8+Ky/9/OGaBigiNYQqY
wQ/V+1IZaH6hKDcZSQYF7O2HJajLCmmLZf1dFxIv638zhouwqmjN6JHJbR+a6RlM
olyno6LRfngXfF6RRoUVeOAMatQ+u5pfzBUtYUw+gYIHrID/q2f1NqIX+Fr6dW+v
bYnYxtHsn+ICBPs1Te3eXsr9331zjT5wTi5RlLHxV1wKZ5i6fPiFnrEqPHPGtUrA
4hTBfZ6ICkRO4m0Zzl0zKw5cayh6B3d2UJbBORR53uKC/9kY+hdZYoiNCvzYI9Vc
C1mfYen00rUpG7MmMoVs+yhzbTUIJ/IFvRh8LbiU8bnpc8NeNw5cRj5PjgOVmyc1
XozFEENHSlD7oleyWVAAhOQaZZY9Trp0l0gWU3+mas1ODFQOZ9oLHBKuRzF2d34/
hzuwrpduWLjF4hwL5d9n77y0Aewb3uYK7JoawwMsca+/oA8i+1/X5g5UUCF4LH35
kdKZj0IYfzV7PtxvR5sla8w1/SQ/ElWV3TO5zcJQQnTq+cAh9NVgNO7r2a8hCXu3
R/CQ7jRcOHjov0t2yEbwO8gzsMny2+7QCKOzQGICZWQ6ZhI/6suur9Q0vIrpoM8G
7POfOQbfd9ls4RFTgMgbcSGNlOAU6lqr7o2RWhWgXsgtJ/SdAdq36URhS5tMu93L
DieWkMO17jm3kQgFp6A/k5CUSl/s2Lf4k/suUzM5ScZXFBHOsHYhmhvzQ2uIF1J9
YbQQGnypqD1Zqt3MrRkPjKHnc+McN7tZrl+K0J4xPDukFAYGSMKyNPj/xlDzhWuw
W+ANstKlKSDUnyfzsuETKdQxLnrOUBnwhAO5OdFsLqdmOhIRa3tUpZD9ZE3Gj4j9
jyJCwbMnpJnx5PglfjFQR/3YvhMkQpgElwOhMFQqCAsR5t8IkwsW1kAFdKVo7c27
fjxlJehtyyCH+MDY1h3wkO7Mfy8yyMDVLH+Ut43ungyCizcTA0WRWIFePhE4JEPL
ePEhziqnUMb0SpBCgKXLwxjn8DwfeBBwmL+U/BwEjXi0md810GyE0NB4V68g95eR
bMLw+5qK2kqiC6KhPdrsZegdK4qeZ7QcpriFm5I/aVQ7ETpC3Fb4EwQZmnSdunc4
/SwFTTU7N9MTM1hNTk6RoXaU3dmYzo/68x/2Qou4bjzVxPTB39cPB2y1N9d4QxsF
fW4FOBz1zNjd+MdIO3QS+SvoACkorGEs/e3Z6LfDAoKGaq/xzNXvRf5suIH7BMKT
DXP9rQdQOaz/otB/fEAbMG5vhy4ZZhRu1FY9dv80JGy7dSd79t1a95vGTMDxNUTw
KbaFqUV5TVDBjhTdYvzKIyOooQlPzMyawXSL/+41G8tO6azxh/pRG7Xs+GXvwAeU
F3451ja7uy4RrFy1RkGCuSu8Uezcd6yH9RmXTcp3FVrgjUmS/aX7+gB1pCIW6fR6
nek+L5Mp0jdpztz4NHe+La7ARPQuuUxohrEwgcTWW80B98knMYypacj5Gi7ywPlh
FT3NoL0xhz5QjxWMEk3Z6Y4wDvO6b2eLdGlbBtBE5NUXAzqPi2c/PGaxt5KA8fFn
p0iKsXrb+5VUxdrTAQik2Uhir9/EUdfJLblZWjRFuiT6lyodMtF4PmRrY8l+v8f8
1dpvj9+KiN+UMtZ2F6MAWCqLo0BPFj2TYikoaM8b8WTyAEM97kSsAFLso6PuQIhy
gmZdulIjv3DRose128X6NkbH4RqlAqhaXCN6Pi8o26YYNDnlRhDtcJRjPVSJqy9n
WFe+eugTxtStxPZoc+IB6ATwY0cJp21yskOwcySXBykwyodx9I+45jOEAGJyMQMW
HWlROijmZ1wAzV2S+48p9JahS1CvXEdLdqMRB+OwnjgChSeUkNcgvDylOg3EhKrq
HZqTLajoWb01GcDFKFVWobU81F8vw3UgH7duhV8UFGJLNMtlVq1Ck3mUxe7W+Col
3Jzy2gbfR6Z6yO6HilAZFD/MTcstoXZPqeJDs8ibDCr4N5FIvUvbGjHzFF18G4kA
VqnDG4X53YCX6rmKwKBlyG648FL3lPom7v5wX1F+qgzayLd3U2czWzEcntLfydt9
3LYWuNAkCHZWw4vfqSRTDavgcanJWZmD+38XAEH7FhKCezpHECXuVqSVVT/axYKz
XQzAKHLIMx69vxOWXYvPCr5RWsoVI0LgXKrqCyg82bSwv2C2K+g7zKevD4ywxqra
Ftt6WE4wQlypik0uKab5vU/bxgCf8qtIMjujhZcNq3X1oMvyU76joISS2eOJeqq3
4mVNqiTfiu7NMZMbWWRBmUUWtDnX6h+96pdf7APR8fhD3f4c03Sgpiaz1XWhfISP
J5eKLc3BCYS0TOjN4TQpf9pew89+jBueaqnHYh3hBCuTLbZqpNT1OTAd2bWosgn2
LMijA3zuQN7QuYOhtHUkQiB/Xb4Yx1L8rxF06zXo35qLuqibGL4w45Y/FQqfZehk
8THINyZkezrY2qG0qSNUA79OrJDzDbOHuQlbwyU9+vbIkPXJmvp6Eu3Pjf0MWgjU
l+BoqiuNSgc4UgYWIpsZOmfJib4r8vyChr0WgSKXKRBX2Zp8u6AAyfCZ4rk5lhhl
vdVwrP9F3HhDSau/XgjkIpR7PRinEj5x++ZHWid4uMee0Ak60pbE+p5kxDB8JP6p
HhUB1uAiiKZFJ+kVEWSsbTXLD3EtX0WI98qmvUhUALDofhaqWhnRE9W3bre8cjuU
6pkRaVDXu6RaWFYGVF2fIjou7ZwTkzpYYVYKwRroqfvSZk0bsuMCjfS9bLCZUj7t
y3tFMhkI8FrgKhztGzMpuKS+cPIHHk5/9n7cQSp4s37ebwDqSRDNzF6sDnQ0vSFW
1nvlwfsLaZCbLx8jRSVWLqudNIGEyInbXkotoBdiVWv7sdYzIvk/RmgqVydO31Lg
Dm73m5FZYUij054BsxsdW5avNVHKx3eo0AtfOwk0exA+lC7D+bODvv5dsvRcp9IO
+3gpP6oxHx9WLsLq/ximpyNyET8vZExJjuLQK7KQh5sO5vl/pquMqN1FajYI+HFh
gKTKiNEmxEQKmMBzSLDP/XvKQN7vubpj+WXedk3R3f0EHDw03qr0GAAm+qN+eTyo
ul03TIg67wQ/Jr7zEg6MXx5msEuztLqG7SZrCuZ4C8rpHhuRN4dAGT8oapGvZfGH
WJcNsqFT6WnQe+gIvT96blBZy+GhZ5AybKJgD4/K+iSzYj23fu0rhbxJ1oKx0xy7
cSAvPEQ0rUBqe4PJhLQfAIfUhk8Ro44o32OACohKLCG7CTb1CV6cwFMmnP+4VV3l
EhNevLY8OEwB7DObjzA7sFCUpx/GdiK0s/K7UuO5Tb59kP70B17oGu5389cDhkeO
7Y5U7O+xBfvBcSuy7LhdbCIWdSg7ft3CqTTU89sySPlB7qSOiyM/N2TJZRxMlidN
rdx5PKb5DCPHGfrcuso1IuIsnxAAU7FWTmmsq+Dt6WIqmsn1ng0RpmIWIp3obelb
p6kQajGH24UHsSKcg48qbJbon/D0IJHj0lU3bQGY9cWCtefSmlepXJCs9Pmknzbr
6gc2ctrO1yvH/JqEBm5vXXk1CCWuBpRm4WkqulCjMJRJM6yMzTSEHN9655SviGz/
gH8FkHgucD/9BuS8qGef3uG1ZPhbhwuciKsF75Qd4W2lSZUxKjBmux/TQ0SRxgIV
dGIz3eRdajspsNn04z8LYZ3oeIQKfsCIIP33CtdSfT0xocBKpTT0PaIajxSy5sEu
qGGXfkW1MNdR2xmISN/eHtSdVBgSS629qUHK6N4jb5PHR1o88djOIjfOC2vLEBq8
4Ls2MBZxByohJUtZZEX829F9JyDV2Co+OFtnpA1gcQRW9xKX9jX+Am3TvrCJsOgu
65ZjW3RGJddEphSqT/4Ed2cFl4A7kDIv2asRDFIQcG55FDljDw7Haxdi1QeCztjN
nHIGozIHsFEbifOZ9AgTBaeGzSfMAoriHNloxoqk0Jr0ZmyA5oHEOHD+bjV+Ss1F
2U5MO7C8rkikw6scW1SmSNfcIY9kSPtXD70zJ2nTV77qcmxJgNZnTrRDmbi2H/aR
n660f1n/8QYo73hezwHHzOoSCdYww6/AtLu3M7t3/NkkiaMDXQ0nn//DMkbd9tpP
VoncoMjzzL2Wvs1J9irs1MhQCwI1L0D5C9tSTjf8eQYvpQY3ht7naPd65L8vKJ4l
Ch6bEoe2/15YFuLQ43gD2Z/+otEf5Jlhrm64bPlZUXCUr0P8shmccZ6ccWBoP8wW
lPIjs1c/y09QLlrumQi9n+EkuyGVlAl1ubI2RV/zPEDyHNHAk2RGSYLP4QcfHkKg
M9qy4ylXSqzXLTetsq4bY+KxRHqC1iBAUMAg+TbBwut+TjGLqxCtsT7COGJCxuDz
OVK/OJ8mQTsY/oZG/WmVJOuE6aG2HouyLhyn7UaksWgKaji0CaW8En6wUvflY9FZ
ZeK2VakjCBH3/k+gxa8CAJbKqmPCW4o/Nug0FkpzPoGpPVyhqoeVfHrk5ExMIcXu
JDzDulzO4JrAUt51ErkkCUnit/Bpanvnil2YmU6ODmp8FiSVgdY2J3rwJjI5qlep
dWmcVnpmhCDrJrmGiKLzjoNTab8ORflRgxHnMq+9in7ydE40T9JEFhYWmjK+f1g4
MakHIDke4VJY6X3TdnF9zl5CZ1gjLeinIgccBlYTcWGr/NIuJaiqXdWLdQYRpRzu
7zthh5FWIddAQJOUD9kldTfYMkC2cQL9Z6lMKXqz+xckyg4bvpmdI9AtG2P6Mr4M
DIfgtNdop0OUMkYj8s/Dq3wDpiOnvuuuJJco09kZ0Obs1K8Y3f/cvvtejB1fc7CE
t/2vXz0VxGCI9m5FV42DjqlFV1wbvruBpBHPQ++aEC4wlwJiasrc9gUfcKWI/W0b
2coXBCtXuDL6RP3+wM+XOmkgddGON1cGgjIa3UmrhoYuGNKusFODCGmhvnDYy6IO
lMptCNVfeQKORXJ8eJpox1Sot9ZhOMEksiUpI2iWXyL9jxqq877Pfi/wPJGsDnla
rIDBTFIyCjTajBISDO8chAXHuaX9woUnWUAjkmZ4kCc9Y+Ln3a8ny9sfJieJ6LSg
yV9PolQuuaTlVUkSCjXnYIAVy10arUt6RfQn62cRVM04oobP0WodBRCEoblTW6fp
i73xo28n0yzsBfI+CmWNm6bvV11Gic/cY/YcoWvmohf5U43IdtnMAY2RDNRCiGBP
pRwXAfyzhL3UjPgoMilwGsmxGykP2di3rxCYIH5FUtJ3FOMgc6q0XRiXEyiy0AIn
tTY6L+zVNlWZTncfZFAt01he5TAtu1hkKVp1VsaZvNHbkuxe8ame0Z27Ra8LTv5n
jYkWs+2sEjg/kbuFVDg6ssFw9+ZjCLCNG91R041hzV5n7DkXZMjsbzXpwaaBdtf4
kZ7toL2+HFDofq590MyCJ+U/ZhXdWC341CWAMVlNOnAMm6s9WGF4EpY5INuZNbCa
ifBHErokRVJjgvYoSk5BbpxUmlU0Uxhtb9e20mie8wOewrD7dFnnu8MlqEQFb6pY
V+YymIRTnBtHP1B/mopTNEeqr8M7yOtCAVN5GUe24C4MH6Q3HbOHGvk1Gp9qGw+V
DOJZwTlbKii51VFcPdNWDukyzOmAOvdfpMehG2LuEKFOAH9sO2Leac9mJTN1AeXH
RoBW7hCF3Zik9YJtFFbUw+CVpBJP0aUAzBJQJ0hAbKoybYaeSl+EaTBNGvxdEk6y
VA9pVPHpT3kehWTejsQGIqMGurrSo+sVArIfzh7OjEaXRxJj0J1BHx/vF1ZY/3Cl
RObwiOKGx97XpX3hYWbaljGQ6ipN6ehjzMt1OvzPzD/kJ+m/BbMQp9X9rv8BOOkX
BPbWv1sMgYwAxvKkAXVJUDtK9kGfJIxUbyspiD3V0UzsqLLEa3Fj/d/txTcU0O8e
9nPPkTIQbiQTXJxrravLwe8lPZ2Nyt1BCeT217w4htNICENkKzqcB3+CRF8mqcyQ
9LrIAbyqXwtGHJJzzP8hkTeauQzClmZ1JWZ9BktYEsy4bYC+25ND1h5ouCdfxWbq
vLiur9W5q+vpWiyzVl4XcMtcilS7Hi6iMA8WOHWDe+Sx1KHOzczMCm2W0nZiwh/G
Z73gpf1jI6TCCcuZZr6a1yU9xzC60PEAb/pL7oXbHcKoeyRjKpgPDifrX65efRcW
Yccc8LCa4snAym94c5AJ+UY+G2s0n1QMuXpojnlijPimmMSYZ/6X/eDPEZk8g3Vh
gBCgMCM5hhGA2I1ojw4hz6BRNI2KcGGVnrKm4NOnZ8T4yBI/dAi3RG2MWu7vPch8
OQyF7acsR8Umf3Wf7Yv/KA42E4lSy/bUiOOSN3p+VTs4gRaCRJk37XDxQO7Cc1ib
MRIIhukziIeXBg7bxJPlv5/brV88EHY6HGVheHreT4cTKYB6NUHvp993Zq8ml5Bf
bI3dVNbTqCri7lYjnDFUOxFxA380Fyujh030QNxZlmIfdTLN3zgfdjH2v2cAMUhh
0NQ1P+QbeKwjbeLLEArYTfq1gX0HfbbEnuaof/xGlykq0CYIm03sCiUf3onky2e1
ZPI0QqUEVXjv/q8LiELfCpAzzJ2TPEaDNUqxx0ZGlTaLl4FOsWyyogaycaLYGkPU
M1fD337+BZmwEcUsw77etl7cbSIIkUdEnoDKe3Q7MvialZ6HZolFeSYYmfOBdPj3
EXpgNgs+HZkeZ5apW4o+sgxc4/+6D+gusQqpFTxzaMEFBqRbynnGAltethgZben1
Mdm/D4z2T3iWY40EmbOg1rsTfMxspHB1SyxacZ0rZyoJqPz8LnX3er83aTD5MAmG
D9+1UjSzTfij52Kk+cgdLVG73bdOCeCPQt7mDU/f9rnhJY0IDsUsR2tgMNdYgVLd
2ns5a8MJ14DEf6R8CHOIw8unh4Wl19h22dSzq+Rwku6mTq039NzXpa/nyHY8exmq
jEir5GG0ThA7stiOL3rNfsIO4Q79JhynHawsde9GOdY4S0JzFpzeEVIwqqGJ3pxu
tOJBjNOHZPljRge1lnIf6X2V2atGrTqJzhNimlm/R3B7MWMsrF6jWHqgVpNvJzPJ
Z8P7MEtfIvAi67CToLaDA6BtRkW6FrwNRuu1NssJ/sqqsnQdx2R4TljFpr9qqN7J
jC0nBRrcacv9oZw34/j+ofqb9H99W2BGubS+/UsaaMukdLkAqaFBZSHrcLMn1s50
L7wUfFKtsSCuLXOJtbSCaBJ54TuPzXIn2C8lIlMpfKx3IlcT5sTcSnoOsuoljJTU
iuOfsNeOx2OJrRQLt4gZu8mfX7P8BHGYhvQsWeqZMhvuhLwJ45pszM/Wecn48Lho
QoGuq9R3bvKuGpEILysDmOUNMOE7rfMKkaXxTa+iZLaSI2aiZI9ZKlKczKlHKL2K
TCDZdrbJnoq/Kj5u0fgtWWYofi37x5tV0e8VaQS2LpQNh/W7kdNQfH70d8b3f5L+
JrFXN+4CY3ygOncReiLYtTf6kB2uyKphJtpGfpZaaNKOUFjW7qg+aVEyMysEjnuP
eKAMDZ0REUIvxDumH2H/MVvb14T/nlc32HM8kd9JIVYH9oVF9xYxzoI6HFXajUvz
nA3fkxWvT1YUI9tGDDKnEEKNLCOe6Jv6M+DAGF0VC8mwCoLdN9Ec2VW8x7OOx8oR
3LMpVCRjQjmRXPcv3eOHoZEEmppVT+UTu4jgwX2YTvM+bHOw4j2/J3lLchG4NJi0
GuyKXoxd/gKRqllYq7IkurRKVcNvkw/6hIoKKhWTbSAO2x2WyyTDruqPyDN2tlUu
xSYpylhwQbf8rTAUVYe+En33ictV5SebUrnCr5Hosrs8MHOFEbeuY1Yr+GY5dlnM
8eqmuhnVHwBIo0JuMn/CqD3crY9urWdoTha/Y2A6/uCahjM5ywU0eYekw867BR+E
Pz2Ixo/vErEJRjtQ/7EmO/kaAW5fTdUKTWroYalzzRxNoAY/0brYriFyr/D+Tyv9
nQSVw03RNX4UD55I5TdvWd8ZKfuhANlTm1c2zeE5+AwZSFvycoIUyrZUBF48Y4JC
p/1HwrqhRhViZ4wUc6aDznVr78zoTpKMblHkvd8mLw3V6B71KXCy2v0HnTgCpbb9
tdyKCPzFeQ3ygrEP26qqUj2uMgBm9NGMHUnOZ2+Fo0EbYObmKPlSAI41SNTEyu3m
JlIonx+ZYRaVsUu5M1Tfk2xSkFx/BCBtXfIA35e4XMk8D5K95l6b0lkeNX2N0KE9
FIQeSUUIvV9dHbChJfYrb5qm9XtpTAA3EHSHYUR4mMuaFijiNgLc60yYUVxMkq5M
wg3bvqBtQt6AljqUwhuljeCDNvtreRsHSLACv91siA6xq/E/1pWouOwZd3cUuOH6
rGrs9MWvf1JYMuaQHejDAA/dXukb94JGG/pyDtKojvMe2V5ctHv7QaV1N5V1Jd5V
OgWmEsiqIZKjEea96J5nfukyO1swdET7QPZYQhpL3KdQqWsteu6af7Y1THJAbdH6
E/95r00raG4mJcyRssV8x1H69SjCewVQYD0ySI4iRx6IOQ6xZUXrmFYlgD/I1zCs
dumtZAmZUC2OsoO4QB07juj3s7jHyMfEwA4T2dsXwWKEZZuormHnRnUF+5G6BQNS
a/qbxdWmiDQFwp1lQAqT1F/BiuCQls3kN5ss1mMVQOnKzdK/54uoYdkQsESMsrxW
mGBTot4w7jIs1h/OahJ9hzE0amKpqTTQJGsoWTcPDK21TEOu0g9ciYbvBfpnoqe6
5maJi49gMFfLrdhr8RFFN01IIOizJ6xWoRCI5PholAWP8G8jdHWV/KmVzlsd80Nu
wiDSNfxi7qme4Zfy2kGdL7hNBAFfC4kH/sGfchYYmq3wekK6O4TVvAMLKrH3kWmF
/AZjQWOCDCaB77WoikkjSYi3BSaYSJULzrdQWNPxkQicOhRxbCvqfOsz+0Xh33IS
vFvX1yr7PmboiIExUbkiEX/bEHYVmRiWUpQJqb39SXaCiDQ5hCyu1abx741onw0q
HyIp/5z8HtrMCV9iwfKcOjiD3A4gqjEpWxohCs8dzHq7oDJ3IkrN5Amw1e3SEJDw
BVBL+cSfbAn60ttjoNt1yDFwF5wKIGzMxTCTAGngZGHQCFYQmHF9sh6ZiOkT4wMo
x4Q2a+Z0YZnWbAYhfq7uF80iA/f5hgDEGewPXEdnN0DKnH0FE5QegldjZSHvZW9r
VjCE2hfHLxcA7oUPhSklieCEO7myh2SnwWqpD8a6/Jsg7vSGAyMyai8u4iau/r9w
Im+b/z8vblmuovEU6d83lvusv1JxGZlbQI8nmotBehPWvyWMdKUiE4LyGaMJYqi3
y8vyKQfhTZvtma254HgZwz+uBVZNIa7vTVF4cCVxGB3iro6luauzUcwzDxusO6ap
404nHyVpM6T80U2c559iwMb7919H99T62I/UXj1s/E7p7HT6Cu3JQuEKvcC5cfg3
WFQL4vto7eb3nsKkw1LVFL3jWfA6qRteGU5ka5zm8sw5LTE6+IB9Io0iUcJ64kEV
zEdDFyPSIGCsFqNmT39n8XAFNf6i1C1zyUWlelM3+xlAasGLkrLqM+mIxqvOx/8g
e+//MjI6R8X62V4b3mbe/0LhDglX/Pj+hf6vUSvnvQlHC+lEcQ8ZmGFSjq+UHV/y
gHxXr9weTmN56ktFRKBoVaibZyp9kljT1rMuz0Xubn5z4YkG1t5+L6NsCh+6FT21
V1z5BXgttgMQByfqffQPI4TjGL3zphxxcPZydZdGp+rVpVkX2NfANDzmF8za/dkU
HFL4RJnsYGz9yDCu/TgKPnivtBopUdW7jeBYE0B1K+ufcj9nSs8phlRUfo1aRan+
mI9QSsCrJ5J2ywziEZudmqr+iwdK89U8GdUEO4spGJ7WIpZjxVVyAAb9gMgAH5+M
npZLoqWAsBLOYncjrC/WwM8aqIkWcbs6WRvUZZXKDC619B5rJOg3AqLoq3laW+wl
hBfLgsXj/8lpy2OOzaFM80iqkCDtnKxBkMSnSdxnB8iPxUQYFYN4JPXMUwsdHMWa
mkUhWA13PY+J70t8sAOgXdlO523lyS54lvr1gnXMs+QBu4vyQSLQgserqGdiaDkC
1BO02F0F+irpsCfFnuuydZIIwR/BOO8gpPpizWEnXcsh9G4/JP2B9vHtSkL3i8Zb
jUIVN9ldMbj0ygCNJrUjb5JSF+8MQ3vd7M2T1LyGIkV7CjHS3bFEYE3f9LJ4Mf8A
0cb87O6Ku9u91h/2iXag0QTxUdkZJ/QmIS6LdPefcKnrMjqzVU0SvVPjSpmLWz4v
jAQP4irkhSYF4eSeC6xaWlxTlA9kVsMthaL/H81Ma7Hhze5X2NMLPdA+UHDU/TVH
6dwf7OCCbN4gaeGZo4CEX+mvMTRMlP/lm/qwKPMMfObASJ5NHcJgNxJ1HrENhHL4
ox7tyzlReYbvJAT2rpEcV/34mX+Awwdi1n6Z9+tysPLzzqqKgAMbLSOlm7DeHOaK
V0ljxGJy/vOMXfMxeGjzmMbhbUj4XuuMTk6ZUKYfnkfwUlxdNbbn/zoou9cmIYiB
5ouwhjvUE9Bn1C6g7pnfjocUoLahMZBivdzwJBcFmGXfJYhpX+06y2eR4S1vL1mT
zm3O8C2VesIkAajFkaNQwgE2Ah12YBRSQpi3/Gwa6wgQ/ToeduasUGVAR2ZIMNUa
Wj5jvmtL9BJH/+ZekFRSdRiP6szuEoxFtK2taHiUJrI3s17UPG7/CUOORgTyr+U2
5RMM8Wrjg+tDrzqGwdbViaIG3Pa47ZosRg3Q8wD3eOtLdMkwCJxzScRkuXJLi3l0
TeUA4HHe7392s058Bp3It+makC0xC4Wj9ucq8kSEd9MlFQjE9rPNegwcJ9/2s/lY
0qljfZzhfPQE3f1tENAEyRyFc9Y+x4W3ii0hd0CiykVhiDWVwHcc2yPL1dJmpSBO
dNJHUUDxl0ufLhRetdYozqx11YSYiyIylTHoc0KfgVaAKaZ+wFvOlyo10u6A4fJm
MI5pouYTXwPPEAJ98A/isCTmR7igr7DO/qG/m1uF43Cl09ZX94yV6DLs66L7he8N
Zqz5omViJPyi6DeYQpob+nEnwWMxcHlVBC8B3Ut12w4ixWLBSC19GX6ivW1hdBhx
HCl9n5EtqRPWOcZoQhdM0ntROq6BLLx9ptMyuQ8w0rXBWJY6mcRkSZdFBBs8Sr0F
1psDljUezn8Fllu9QuTd+QAdfaeMsYgX7yjMtvGaHe2II3BIoRRScZMoHEcugmEy
bsDELY/WFwGFlgTGZMfHip/l47caRaLF3wgJ5gbEljnuyjNPWs4YiuHqkKLsVjrR
U3AB0jXtvxhST85VLpJyypJanvWFtx3zyHWn251A2t13LTxfNWXqlj6uEX4cdfPW
2DsJ3RBc4H7WNuyW34JZNDykPBbXuz+xw/KMIEUxrF27/ke3V/EkOlEok0X5YYOS
yBwlEJvSjnZ/cwzh9dsJFQ4+lfVrsGtUAOlhGdz5fGJmJHSApHJDk1rl00J0rodx
Vj8vXARgNUpyqn1LTAVG6BJxmdG5SJOYMOK11ZYBuAHwyUctUREs0JBi2VizKXfh
6oaRLNm2eR6yw140rDY5b94697QCR2gSDr7a79u710vLR7SIkHmFofy28ANXHOKi
f6qlbSv7gRadSiKLhCd3NJVgnCJYVQBEVDGj6aMbbNsMLJqqj5P7V/QH2lm76a/D
a+oI10frXgvBXzUDaWq4/rEOIBwpFH544QlwllJfF/qiozloLWJPeZgoOG9NSdur
/Lt8mneZtvPX/EkUKae1feDAbbu52NtU7125RBJGs+KE/Oq2UUvkDbvfM/nNtpBU
HXuVVoGRRBHVeAti1TDj18h9dItgpxos1YIpZeYPZUrwKrWvKPjC73LXFDpyzPSy
LaiUJx9K1Mgf90MuFlg1gCZRVICl+rQqw9xQ7LB3NBsogBrZTeyKg7bHFXrvVT3H
rajQjkj9ikDQzcLVRrJxpGxMz743LfO8HqTytcGRkq1RkVtuVqny1xxo/elcpCxH
0Rfy29kimE97xWMlm+xnRLciBqpqTSNd4caFH6DiF0Xt2IFW9bDzeMCLh6zWQt3z
LMqozIC6l0ILH/f318d1ZPGkC6RVlEucc91VPV228ErNwORlY4spvrBG7bCtlI/y
Cbj1t51e8vI+kfVCEwHs5CNSLoBGZP6acZ6GkIm3eBWKehSb58G2aBhyqqWIrtJc
sbcql5pnmXcOfYatkF6PlLP/GmAOYin2YJN3kMgBECPQdp6QqzLd1M3tjFesboM7
2j4gS7KOQxM5yp7eFG53A9m2ZF1mR0O4LaPQo7hrhcsRNmrFEYkXk4cRck32Jjo4
jMu0B/2SPfJo79nhS89LW+263GZ+ttZ6dwnrxbYhhObVqyqB3sexTrIhjhSUd4aq
wpDIe4Fs1xQySOyuLb1E218um9P+t2+vl3co1ds2z1FDPmmr0W6xmO8SszR+CxUQ
lR+Vv86W4yi7BFde/IH9sp1nVi5OCecj8daE7ygabkZ8x06VVYc6vMWf2I+S7e8G
to0JRptLhPgLxSmQndJZs0NLhz10al30tCR7J4ZjI0ilOD9NhWuu22mDvV6kTobS
Zhd/6Gy9BXrIePcBSkRGPTIs4kG/Ppw6VSWOxR9JQERenAxIaNl3Ro3PY9eQ1NmA
MGEa7N62NQNd77DuRe+53jbSIMeBHvqXft+R/nuFxVIaKC46fdqAeFiOGzdbAuC+
cA/yeeNvNknL7QXhJeUSN4f3C6HcDDHxxu30UJhr1FzE6gTfv69Ko9HcdKshBwHi
tki+M+oX/e1qq9yZHq73XIHhZIz4l9sI+MbUXvANsjU2iBjoodLupGz6nqQIYwpH
sXQpld1j26eycVa5Gxsfx7KjIjFjvT9tAklUOoLzTXCOa9Ky3o5Ad8HuuUmZX4Ed
cXjKSe9+zL+JfM/VyI9xQ+0eGgaV4Xkt/4PtVMIKICf+PYjpVaiwvRSLT5CqS5ha
Wyy26ebWOQNbUkV4IqBaBESV4zHeIty4rrM/ARJ8UMrifTukCdS7GerL8dGIARUb
wmw4CFbUx+kdQKVPdHM5/04DAgoEYSX4Qu+AQSrkkFfCLo+TQ9oApjUrGYx5SuCz
Ffh6aRw6DnvambdEwXxgdKJ3blT7relC5ifdpzIJzU9L3r0qrkciLlufsV2pDLD3
M//qkfgBQV8bw4Rafz1TlWHIPR3OiqxoEKZsVraTVrr0D/clNMe2hmthhTXobH+C
oSZEBfGQLe/p439PGambxP0rFc2Nwlze5is5dCb1VZsVeZi1zvM6Sq/t8GcqIzgl
ka1P1O7Dt3MLf6B2eVB9cj6FCow+81Us2rjgbnqAajNR4X8ErmcMjMqpgcgSnvmI
7evEp+Jazln/xyo1rHO0fvZDxN4yvsFe4PslZ1oV6s1C2SFHUFp+aqgAZDGa1WPq
bU8BbhARgHMPPsMnp1nX7pkVYueaFF/4MnmFAxlzbkE7TbdJoINPtC/X786z7T3C
PdI0Fm0xv+Iet9C+23aMfM7BiDTh+Q0UEtfz12w/9YtQ0IEtrgkZOso+SMeszDHQ
1FS38M+BcFIKqMo1HBKN9H8EM5a3QJC748Ep4ehPanBhX+vX9Ie+94WgnNsLZk0Q
mU0xQ5HEa3sh6ivkey5R1IsnF+uWLpXSky5GavgP34OhaSegjwNQwtJgDlxJhekY
Ef1CYN93kH/Gg2Rma0J6ww0Fl1rWYo9Uv02PTYTnvxravZrbMUPvRRHXUTQnE/a5
qzZwuZN4ZBAz83bCeRzPCRB86bVuTmwqYeLWV7KQmaAu4mYujmbu0gZpED9Knhgg
Zd455I++NDeIgB9N7vMR73Ew1ngdw8Kxn0YDf8bDSJK6rcu+2Fvh2rcFNGrQ+A4f
cBTNhfhSVQAxvuM+OS84OAAG9UVzC/eZT9gkS3hnRttepGxFr8CPfW/+bMuwUNdj
KnveKBOnpWMeJnSAkdS07XWfVLF7y6Toz3evzR/aKoyqTlc6+OyuO3EojNbpSNoe
CppV6pxHLFmC93S43C/7TTxm/iWZAAu5t9o01H5soqohhXoybix1t54EetBhwtkf
qzXPVJpeh1yyGealswI1u/NoeqIRGeWDcZBgdeGXZLslEiEMNl2l4ixHeprC0FDW
oWX9JeVODUpnaXQfZDxZqbquswtDZ6zCc55OUxzRpjHzFuKjVKh8Wntt2mhYid8e
4qj9lV6iM0AJ+WgbQ9TWgwPUfOzhWIMI2DKG25jEHcMJmNgRScZAksk9IvThR5TN
TSmeu++Setgga/SCWvp5s9Um2NM11lZyxN23sdbgYQYlZsh2CJfvl8+opILvZthv
S8wNHv+BLynUlU/tBAIPh6gM04j/d2Ka0Su3w16xf0Ies2KTI3EAxhIz7Kg9U+hf
Fz5qlmSp5bzC2LlmTxK/IKUGNWzgVzq0Tjwt1YltB/92npRjHi+XAPix7y5Sn6OA
+Gbv2mD1peDzScE4YXFBKqUDRF1jrCci+t6ZQz3lzJsG5H6zSNX8L70/do8oZofx
GxUlGju0TQj4kIeDN2XAxhPYBjz9MaauMHEEYrkZ2PoGwEy7ZsD8Og0usUOLVhue
eq//F145brXqmnI7nZ0nLFOLWanbL32OTRtTQePzkWP2MAmT2DY4dyRTacyZzeYb
r4xeKeubcNOf9f/jgjqn7kFARzU5pXAnmn5Btbj6JqXhhzbvrOq3cK0l8jJLdrNQ
IBBbf6nXWZi5YyuiJIb6wc0M3jl65ecMh37EebTygUUjaYUWHgDKannE+GWO6GYK
MbDvRBNQhfoVkKKxIAW9cF53HyUXeaCC42jcAHim3q8bsf+Vl3jHByCuPwuXNJy2
OKub1z06CvXhKYue/qJnLnMfG5vWViVuJpAKZFqVYQW/JGCyM8sHCbV81dmyS2Ae
0WKqM7M37CYdXXFyLDYcMzWzfyP5PAMslOdRvU3ReQNPTfmHarmPjAVIj7ItxCxf
IxvlmFH384Yowd9R80G1SwOoUnaOKyr+YUZRboSb0DgcG9gsAkVrCoYpJY/inlOj
40eDmxbi8+HeaPQucGXQtr/80NPVf5q/0OhyMJZ65KTzvFCuIAremShN6DbarH4E
LdUyAXxTS/0Vt1llShCyEFjVf6XcXw/D6dLnEStlOnK5/EC2/SPYSByUgj7OzlWn
7yEGMUIjvF5fBMBiw5b4+MX5OPMGqZqef232xRDhf+kngWARo5Dx9VJCtprZ5iim
noBBKMcFc+tOfanX4oL4cwrQSDHiOg4LjrVoG7PlVJoOVoEBa+V7DDbfXtPFpkO8
pC0813F/fwtQOmfKw8lYDEPXw5sI05P5pkDm+1a87IH083DlwneuP4CxkE2l+iJQ
JEuEXm8YeTSvVZt6rM5VP7et/727WXKVIU4fdY/prCYgAXVFDdDi0pKQKye/AOfE
UDtjdGgOppozV0YQLyDi9ZcGS4uI1FRCL7Y0qfjSqPbeinpQ1bx9YawLGXHWrBGn
CEuWwR+qmRrrZozKzrIb03rCbpMte/JWqFgwe9jESAt+UZoZ5RmxLX1Gq1p/vB1C
T8wfZjC1Omiy0JwUIlmKtff24SP7o9L34ziLe3fESfV2h6KA4khPlU30U+nfg9pI
GuGXerouK5mobO3gKpgvkKp1r6ODbvdW2PiZ9if1PSdTGoHY7xK25nCV3DpmBL8j
j3sWfUY/BrSynOJXjr2sd4GOJaP9A3KMxUhkufCS2F5Jcsgsok6+yuSXTVvokf1D
QR/05fEg4WhJpk3Bq8WQqp0XLtMYkq3YSBQRVjwIA0nZn8lPfvuYN+bxiSXS2+bA
Q6SAIM7pLC4mtDhZ3Sz2aAx5uTQHS8KRoMY/asNAGfd2pyryDL9eSdLfJzR2bYP7
d1idErTQlrAlYWITVHXiXRD5ialDjwbBSCWnrJNHCqhQpQRDRe4MaeBn9zCj0cdN
rdcTaYIRHHHSEO4U/2b1/mNd5c09MZMQucwy+c75NIr1ofZv9Hb5q2E8L4GEcfY+
XmS+1vKboipI2zC2OZ0PGLxDjbz5Z3B9wDTX2UqI6QKML4gsP9/3JaisFp4705C0
JZ4TtqTTsa9yGeRwwxt7ISrdeDTZg2HHT6oeOo93uLmhuWIdAGazblmJ2+uQZ3eP
A29RGpWXVw6wV0RIfBPZyWlZ4v3enqkITEQoQjUJEN2vpXMzHu3FiPeI4vXYBHRs
g2dM7qSm7ul+maYRkKN4ybvHhg9nI07/TJJ/eRAh0/190B8g6I8YqF3LWcEFA36o
ovwZ+3mDDi20NmNgJy3WARhLEJXKb8dozbjyESn66CQJ24/yCjkbwX2Sv7WgO8l0
7OQ9z3RESWv529+zwiwW+WOJH3RQhvNy0oHfvB2M68Jh3ELHl7E4geQTuho6EtJ0
AfAwMLJnu4CfdE9iZyP5iM6njXUl6doEMdxB7bKODNaw88ppmkZq0zSA7TKwSlMo
510zXf/Zqnwj+5e8+Y0sRJGm6n1PjPtAdMGSTUmWuY+5/edj2PDGqKanAtRv9SDP
fL/WphLxDmIszO9ikypK+D3cLhQ2eiu2pvUM2sbAcsi0nu5n/c7dv7b6l302XO5h
GpHmd7jaeFV9J13pZ92bUkUfkFpwYrsoeuY/EWPNYesZ19DGb6TfX7+McWKHs2Dn
2qBbJ2NCzhj/Y2SSYT60+1jYngbevm3LYZ2LhJKcUWNWzaZt0kiqM+FwqoF4oKYD
8fb+TdK7pEcv+GV66Y1EAu0JDqaJmpLw58zaRLLCmosDw2WKbSGIT/CFW0pVbEEP
ie0SocPpfPrX74Csy2nMSqx8uuPjXnIr+b4qiMZ5hJVWxJU4ylo5slItN4Vm7/aM
LHBgDdfzfU0viMkFFl9vtjpv0qgHdUe/GuVS6QHCiVkKl/TgNOwyb7Y7F8MWVRMs
qctYaWbwHTAbWj6Uz5Xv7AjAAEIo3mWId5HjX/C/T3YyBK0EkV+pbusFv7R4xBEl
eNPYNgAsFtcg7yLiIO2oVC+aEn7cpXlEAA2KIHznJy0O/ECoqdFNYb+1Y6/pZYlx
TF2dQw8UyZFSLmVGpmB4UV3wr1wzK9FCCeuzYcnFvJZjYpjJDDpq8oy9PFY0tP8I
ncQStz6yXyC0Emhk+PCwUpnQbufCEKd85BUEeTq/m6aifwzygkJTrkcwwUFmwPII
wppbXJYl3vANk3oL6AOnCt/Hlb0YIcwgdq0HuvsVMpC0YT51gNa7mKtTgtvRmoDe
x3GwZWlC6pWr0XYVaQs474zhvfXZmGrlOt0Nov2zIPcZQfq436HxhLzephy4VQu5
hTpsPxTenwT5USkh9SHvnBgfjd5cGdn3WyuZFK/tKjhpolt3b6WodGAQDwFU5Ysg
k2Yn8Oxz7mIHXJVK5S8YrdkACXtCva+hXvzBi/nWEtHU+j0DWdFLeUwsj6HFGR23
GnUBFbm7uDP2zdmpvcOgcvlL3lyeAJfAZHDveaeAPxk5rOAR9klZ43A9KN3CnYFd
UQgB+J430n2TLfTt6f57UpuHJ44P5ZfMZa7JJR/8w1uzIbet2qjaXQOZxsiYeu13
EVUY9ffLqYGUmVBbzEWGeM8BOzbQ2awz5sfWQFlwFLr8J7vF5Cg6rnOtDLjEIbyj
ageawSIw42W/PkMvTiFBNp2A1Qc2H8hFYnU6/7cHGWDwHicKiQjuZpguE8m/JNKT
80z8v9AyybxDliH9iTfKacVoVuaqtrMLfHLXs/qVv8wdAGq+iGtYRYChWTk4KLZi
+DQuSO82PPmL7a/UPlVbmkdeR1XyDPGhv4OnUJXp/e/EpS7knMhY1883MJcuAELq
EYlLiAdie+BnJNdyAGtbb2A1yuXNwEDqzaKCkVfmXKprH0m/y2qtI9CKUeXkNL9n
4kcMgEsNAqYouwOGQPws4rAIsw4tmOVJWAe6rzYZuLI0rFajmnuVy4t5XELmvxG+
qHfau8X+Q1zjcuCccsLwvNS9rCRRO6xuDPXfg0T8vz909LIWA9t9K7nT1BofOf7U
WlJVvHImvxaS8EMEVE9Gkop0b/SYx/JXanrk0qFlakmCb8rDRuYzcFzHR4Gqqh5+
hI00fdapVhEdNK78N/LHclRvNoOwn0SODxHcHQrxCVx6ExCeqWwn8LreSrZp2XVJ
6BjWFuKTmrAE8cJu0FMQ0VaaiTFD1uKhsY9JKsu+rdnOOuV6a1RQSgvoACi7Lvzv
FB2bEd88f9OX8+72yQ88o4nvG2zzTFC6a48NUGO3efWsIcuYksz5jgWiUDBpx0lG
Unga7CauSXxsPfXivkmHttg3p+qDLnSR3L2a7N/drXYWMQ0z/WlJCxYJ0HbpR6Xm
9RP2Fxk1WZE/epONOnE0LgcZToKskBepVA/hHViAjd6tfo9aEiZjQkjPc4JkVpAS
egy2LpJeQM17kkoP5QzbPN5NurxsVafwkLFVqpjW3stDdJQIvR9kUkuXYQOBu/mP
nDhKo76j3c0UpuJpSnj9MDvLLDniKGlu2a1Pq3vkXFNCpLTAH2MTHP/8ByUGlfx9
XLtaaxNVQVdhiRLUZz/SZcUEH81rG4zqEm9EfWB8zYovrshrCTCFukD0kF7fAa4S
tWO6emK6rwaUhtPLHHXoJvPes1j8lguCaqH2gtUuOAcvXtk5DSU3bfrnMb4mpnyT
V8msZ+wPruY/fShA9+nRc7vuk376O4q+/oHymdRD6j1vekWj3Tf1FX9mSY7NXavc
PMLskD/samZHC4ZPl5joQeBWAq5I6p6WJWynFPdbA7pjYN8gK/B0UPn+xnSlbE4T
SRXMdsFI5BFnVaGKPR4Vl/EBgshxQWVwtw2i5FSHnCOWoPdT7NDiHyyFwmQX7//6
YXxDnft+eNAKo4nerP0gz/cDqfCf17iajrIOfXQr4sGcCT/ltNTaFpRE4n/9VaOQ
F2FuPjM1XS+FGNd6qkXH+XnGcypjwerLI7c6efUBlmbF5YEAS7IUSIN0wNa92ZRF
qpp3BVLCTKWzN40Ek2UACXJIZ7PTEiu1PKlj7LzaEQKaSPlwwMPavp4Tc+I9VGI3
/MEVUVXtjG5GBapsTE3LE/8r3/fTqsNhfN7OxOiGAoB4Wgx/D3kXbKGGQGg+IU5g
c+9fFppMQ+4QPgDwq9hwiVpHjG4+PL6/VM/PpOc7zWxIZPnloEKcqvvDDrKYqA4m
NK3aScfNCNo+54HRxfukOzYRClhvGL5kZaVpF0HwYVmuBZBj2wPsFNeM2CCe6rrD
XkaXMuC9QBl86/k3PccgBdiKd34G6bcyG4Pk8WUDTalF05GohBWavfWtxdxTlqlI
2o2SKbT5onbdbaVGqdPMmR57Tdqo58gZMTxPM0ezs3gqXnT2h+4ntiR9e6G8HhMw
FUcVBNcUEtm3GodX21L3BrbSndrSdwudcqrSFMvGsQbdJxbLjt35SGhyLR9dQJn4
5/BZrHiXJHX/mtrk7xvUVKYU654HXalPb/pt2afG5ErACNgsvM3ZDkQhjW5hjMSy
zYgT0XfQXQuN9jq7O1phZMGrmBOQoyO85Uy45EaWmlWg/zU4+CXPyhOsLe7LTsBk
r5EBI51i4z87Gb+//pmze+Y9BdDNUVcOEtzWAvfs9J8ydf9KaF+TIaWv7kbjZuCw
fL1Q97lzwl3IFJzLb63unzrDwXYBT6t89AZw+hkX98WCQXBo8HWq62JvJgmyJxZr
ilNTH/L824jk8+5p1vY8aBWKTbHh+uI5onHe8tCKvZfPWCMPQXNZ6d+sbg6rQBTO
qmgln6msDHh0Loz3l1cW+v8nN8hDb1eAdz6X38Z0M6Q2yWzrsjDQbO7zEChX5sj3
MYJcz7/a6rLx1Ijl3HhfjfrDEBbKSMQb+ED7wXUb38uqGWvzINOtpMPVJ+34EpXT
JVVK5oTSMtdNCZx+N+EDM3GhrOTEXRZdBf/A8AeL3Ti4xpRYeHb9jfs2jFCW6WPZ
Ef4xZNcyK1mVRpygrEzcIs7JSf0AWRmKYOa7mPQeDabK3+msD4nkDhy0hUgSxaYM
jP80R9cGeM8zuMokdiX9x46jwly3deGH3PfNqalEtGhZC2ghK83+dlnSBJ/hDcgc
MUSElJA0GddedJJbbiXq0t4NBO0NKafW6gR13+8mZgQuvEqHqIER7PqVc2s7ezES
9RWRzQWBbdCUKhXWLzZJ9oqCr7NL5xTfRYT/n1ljStbG6We7YwGCHMumVt6/Ucue
idWRyuePzzTBU3Ru+ByO4ZR+UAXMcbQPPcTe7iXyTXBcWSuABbaCp42nxoyGp2T7
K90XDYURRqNouBq+dykT1rPWwVBFa9T/av97JKEI9tScTJCrDzfVVWVGkPoz33Fq
l/pQnDQ7kSMRwu7C3BO3uV22fZQbiSzmdM7gwTDHM1xVrjcPOE431t4K/5WVyNei
YlUnaADhcO1v4yry8Gdet41JeSP9lkWvsSVAX5JO45o139v2JewvydV/plhLsvG5
QOWavqCu7nmtQvjdx/xIdhRYJ4mFyafKMLHgmzYgoQKr0cd+psH+q/UDo3Vt+Ydy
R7/NA7TKqfhrC7BE/A9YBWkqu2e9pJNsZUsDolv/38gHChMX6GkY9W05+3YdQFT6
BgtWwwW+uXQq8c2X4uXUsmnRiw40eehUFtaMOZI2sAk9CztNd0pnWEAmCCd0xJrN
EqQuG/tZl9JY+TRiG0Tfp4Dxrq7gLSQrNqQ0rfZB+EA7FQjmEMSDw/d8vZCRuWGg
JI0blgfe4HaZHGHSxCOkG4TX/zqXIuB3H3xd60EACH7lID3UfdPuJj6UR45u3koQ
6Wc+Fg+wxBxHsV9pMyfCaQAl9x/50fqIQLLCdu8e09SCzHTD2jzCp+qYO7klTGHB
spho+DbcWvcJIpvI1DCgMrF4y3RYZWsHIrao16EozWj8fx1nXjTY66e3NZll5adA
NAFVlUOgdDDomgr1XYVMVMx6w3sbGvvSltYbBY+Qz1ICN5SwwUCrnYKsmSYZh9qq
dTMSaSk3oV4DeZ54lqZdstqug2oyo1UuiC2DhreZMswzJPa2Z8J+S+ekNUD5mFvM
RjAEMq/RdVuiN2ni1PTo5YRTHWk8Pcu+fxsj9bq51H1UDjcEqHX4UINPvkJR/ZwM
9VTHsyUX6p9LagSTcjFnEw==
`pragma protect end_protected
